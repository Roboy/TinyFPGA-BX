// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sat Jun 29 15:06:32 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (pin1_usb_dp, pin2_usb_dn, pin3_clk_16mhz, pin4, pin5, 
            pin6, pin7, pin8, pin9, pin10, pin11, pin12, pin13, 
            pin14_sdo, pin15_sdi, pin16_sck, pin17_ss, pin18, pin19, 
            pin20, pin21, pin22, pin23, pin24) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(1[8:18])
    output pin1_usb_dp /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(2[9:20])
    output pin2_usb_dn /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(3[9:20])
    input pin3_clk_16mhz;   // verilog/TinyFPGA_B.v(4[9:23])
    input pin4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(5[9:13])
    input pin5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:13])
    input pin6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:13])
    output pin7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(8[9:13])
    output pin8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:13])
    output pin9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:13])
    output pin10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    output pin11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output pin12 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    output pin13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    output pin14_sdo /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:18])
    output pin15_sdi /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:18])
    output pin16_sck /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(17[9:18])
    output pin17_ss /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:17])
    output pin18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:14])
    output pin19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:14])
    output pin20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:14])
    output pin21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:14])
    output pin22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:14])
    output pin23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:14])
    output pin24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:14])
    
    wire pin3_clk_16mhz_N /* synthesis is_clock=1, SET_AS_NETWORK=pin3_clk_16mhz_c */ ;   // verilog/TinyFPGA_B.v(4[9:23])
    
    wire GND_net, n14357, n404, n406, n408, n410, n412, n414, 
        n416, n418, n420, n422, n424, n426, n428, n430, n432, 
        n434, n436, n438, n440, n442, n444, n446, n448, n450, 
        n452, n454, n456, n458, n460, n462, n464, n466, n468, 
        n470, n472, n474, n476, n478, n480, n482, n484, n486, 
        n488, n490, n492, n494, n496, n498;
    wire [16:0]Amp25_out1;   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(71[22:32])
    
    wire n14356;
    wire [15:0]Look_Up_Table_out1_1;   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(77[21:41])
    
    wire n14371, n14355, n14363;
    wire [32:0]Error_sub_temp;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(44[22:36])
    wire [36:0]Add_add_temp_adj_2483;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(62[22:34])
    
    wire Saturate_out1_31__N_266, Saturate_out1_31__N_267;
    wire [32:0]Error_sub_temp_adj_2497;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(44[22:36])
    wire [36:0]Add_add_temp_adj_2514;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(62[22:34])
    
    wire Saturate_out1_31__N_266_adj_2417, Saturate_out1_31__N_267_adj_2418, 
        n14362, n19782, n14354, n19765, n14353, n14352, n794, 
        n14349, n14367, n14348, n14347, n14346, n4, n14345, n14361, 
        n14380, n14344, n14343, n14342, n14341, n142, n139, n14379, 
        n14340, n14378, n14377, n14339, n14376, n14338, n14375, 
        n14360, n14322, n14374, n14337, n14336, n14381, n14321, 
        n14335, n14373, n14372, n14369, n14320, n14334, n14333, 
        n14370, n14366, n14368, n14332, n14359, n14364, n14365, 
        n14358, n628, n14331, n14330, n14329, n14328, n14324, 
        n14327, n141, n142_adj_2419, n146, n14326, n793, n794_adj_2420, 
        n141_adj_2421, n142_adj_2422, n146_adj_2423, n14323, n14325, 
        n21486, VCC_net, n793_adj_2424, n794_adj_2425;
    
    GND i4 (.Y(GND_net));
    SB_IO pin1_usb_dp_pad (.PACKAGE_PIN(pin1_usb_dp), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin1_usb_dp_pad.PIN_TYPE = 6'b101001;
    defparam pin1_usb_dp_pad.PULLUP = 1'b0;
    defparam pin1_usb_dp_pad.NEG_TRIGGER = 1'b0;
    defparam pin1_usb_dp_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin2_usb_dn_pad (.PACKAGE_PIN(pin2_usb_dn), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin2_usb_dn_pad.PIN_TYPE = 6'b101001;
    defparam pin2_usb_dn_pad.PULLUP = 1'b0;
    defparam pin2_usb_dn_pad.NEG_TRIGGER = 1'b0;
    defparam pin2_usb_dn_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut (.I0(GND_net), .I1(Error_sub_temp[30]), .I2(GND_net), 
            .I3(GND_net), .O(n141));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16567_2_lut (.I0(Look_Up_Table_out1_1[13]), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n21486));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(49[22:38])
    defparam i16567_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7_4_lut (.I0(n628), .I1(Look_Up_Table_out1_1[15]), .I2(n21486), 
            .I3(GND_net), .O(n139));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(49[22:38])
    defparam i7_4_lut.LUT_INIT = 16'h5a66;
    SB_LUT4 i12417_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[5]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14352));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12417_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12703_3_lut (.I0(n146), .I1(Error_sub_temp[30]), .I2(GND_net), 
            .I3(GND_net), .O(n794_adj_2420));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(49[22:38])
    defparam i12703_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i12424_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[12]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14359));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12424_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12425_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[13]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14360));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12425_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12426_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[14]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14361));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12426_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12427_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[15]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14362));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12427_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12395_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[15]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14330));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12395_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12428_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[16]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14363));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12428_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12396_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[16]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14331));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12396_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_312 (.I0(GND_net), .I1(Error_sub_temp_adj_2497[30]), 
            .I2(GND_net), .I3(GND_net), .O(n141_adj_2421));
    defparam i1_2_lut_adj_312.LUT_INIT = 16'h8888;
    SB_LUT4 i12429_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[17]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14364));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12429_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i1_2_lut_adj_313 (.I0(GND_net), .I1(Error_sub_temp_adj_2497[30]), 
            .I2(GND_net), .I3(GND_net), .O(n793_adj_2424));
    defparam i1_2_lut_adj_313.LUT_INIT = 16'h2222;
    SB_LUT4 i12387_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[7]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14322));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12387_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12430_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[18]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14365));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12430_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12431_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[19]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14366));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12431_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12391_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[11]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14326));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12391_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12392_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[12]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14327));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12392_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12421_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[9]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14356));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12421_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12393_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[13]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14328));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12393_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12422_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[10]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14357));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12422_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12397_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[17]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14332));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12397_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12423_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[11]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14358));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12423_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12398_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[18]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14333));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12398_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12399_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[19]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14334));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12399_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12400_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[20]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14335));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12400_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12401_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[21]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14336));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12401_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12402_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[22]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14337));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12402_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12432_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[20]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14367));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12432_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12385_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[5]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14320));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12385_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12433_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[21]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14368));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12433_3_lut.LUT_INIT = 16'h5454;
    FOC_Current_Control foc (.Phase_Voltage_0({n404, n406, n408, n410, 
            n412, n414, n416, n418, n420, n422, n424, n426, 
            n428, n430, n432, n434}), .pin3_clk_16mhz_N_keep(pin3_clk_16mhz_N), 
            .Phase_Voltage_1({n436, n438, n440, n442, n444, n446, 
            n448, n450, n452, n454, n456, n458, n460, n462, 
            n464, n466}), .Phase_Voltage_2({n468, n470, n472, n474, 
            n476, n478, n480, n482, n484, n486, n488, n490, 
            n492, n494, n496, n498}), .GND_net(GND_net), .\Amp25_out1[14] (Amp25_out1[14]), 
            .\Product_mul_temp[26] (GND_net), .\Look_Up_Table_out1_1[15] (Look_Up_Table_out1_1[15]), 
            .\Look_Up_Table_out1_1[14] (Look_Up_Table_out1_1[14]), .\Look_Up_Table_out1_1[13] (Look_Up_Table_out1_1[13]), 
            .n628(n628), .n142(n142), .n139(n139), .n794(n794), .n4(n4), 
            .n14381(n14381), .\Error_sub_temp[31] (Error_sub_temp_adj_2497[31]), 
            .n14380(n14380), .n14379(n14379), .n14378(n14378), .n14377(n14377), 
            .n14376(n14376), .n14375(n14375), .n14374(n14374), .n14373(n14373), 
            .n14354(n14354), .n14372(n14372), .n14371(n14371), .n14370(n14370), 
            .n14369(n14369), .n14353(n14353), .n14368(n14368), .n14367(n14367), 
            .n14366(n14366), .n14365(n14365), .n14364(n14364), .n14363(n14363), 
            .n14362(n14362), .n14361(n14361), .n14360(n14360), .n14359(n14359), 
            .n14352(n14352), .n14358(n14358), .n146(n146_adj_2423), .n14357(n14357), 
            .n14356(n14356), .n793(n793_adj_2424), .n141(n141_adj_2421), 
            .n794_adj_333(n794_adj_2425), .\Add_add_temp[34] (Add_add_temp_adj_2514[34]), 
            .\Add_add_temp[33] (Add_add_temp_adj_2514[33]), .\Add_add_temp[32] (Add_add_temp_adj_2514[32]), 
            .\Add_add_temp[31] (Add_add_temp_adj_2514[31]), .\Add_add_temp[30] (Add_add_temp_adj_2514[30]), 
            .\Add_add_temp[29] (Add_add_temp_adj_2514[29]), .\Add_add_temp[28] (Add_add_temp_adj_2514[28]), 
            .\Add_add_temp[27] (Add_add_temp_adj_2514[27]), .\Add_add_temp[26] (Add_add_temp_adj_2514[26]), 
            .\Add_add_temp[25] (Add_add_temp_adj_2514[25]), .\Add_add_temp[24] (Add_add_temp_adj_2514[24]), 
            .\Add_add_temp[23] (Add_add_temp_adj_2514[23]), .\Add_add_temp[22] (Add_add_temp_adj_2514[22]), 
            .\Add_add_temp[21] (Add_add_temp_adj_2514[21]), .\Add_add_temp[20] (Add_add_temp_adj_2514[20]), 
            .\Add_add_temp[19] (Add_add_temp_adj_2514[19]), .\Add_add_temp[18] (Add_add_temp_adj_2514[18]), 
            .\Add_add_temp[17] (Add_add_temp_adj_2514[17]), .\Add_add_temp[16] (Add_add_temp_adj_2514[16]), 
            .\Add_add_temp[15] (Add_add_temp_adj_2514[15]), .\Add_add_temp[14] (Add_add_temp_adj_2514[14]), 
            .\Add_add_temp[13] (Add_add_temp_adj_2514[13]), .\Add_add_temp[12] (Add_add_temp_adj_2514[12]), 
            .\Add_add_temp[11] (Add_add_temp_adj_2514[11]), .\Add_add_temp[10] (Add_add_temp_adj_2514[10]), 
            .\Add_add_temp[9] (Add_add_temp_adj_2514[9]), .\Add_add_temp[8] (Add_add_temp_adj_2514[8]), 
            .\Add_add_temp[7] (Add_add_temp_adj_2514[7]), .\Add_add_temp[6] (Add_add_temp_adj_2514[6]), 
            .\Add_add_temp[5] (Add_add_temp_adj_2514[5]), .\Add_add_temp[4] (Add_add_temp_adj_2514[4]), 
            .\Error_sub_temp[30] (Error_sub_temp_adj_2497[30]), .n19765(n19765), 
            .n14355(n14355), .n142_adj_334(n142_adj_2422), .Saturate_out1_31__N_267(Saturate_out1_31__N_267_adj_2418), 
            .Saturate_out1_31__N_266(Saturate_out1_31__N_266_adj_2417), .\Error_sub_temp[31]_adj_335 (Error_sub_temp[31]), 
            .n146_adj_336(n146), .n794_adj_337(n794_adj_2420), .n141_adj_338(n141), 
            .\Error_sub_temp[30]_adj_339 (Error_sub_temp[30]), .n142_adj_340(n142_adj_2419), 
            .n14349(n14349), .n14348(n14348), .n14347(n14347), .n14346(n14346), 
            .n14345(n14345), .n14344(n14344), .n14343(n14343), .n14342(n14342), 
            .n14341(n14341), .n14340(n14340), .n14339(n14339), .n14338(n14338), 
            .n14320(n14320), .n14337(n14337), .n14336(n14336), .n14335(n14335), 
            .n14334(n14334), .n14333(n14333), .n14332(n14332), .n14331(n14331), 
            .n14330(n14330), .n14329(n14329), .\Add_add_temp[34]_adj_341 (Add_add_temp_adj_2483[34]), 
            .\Add_add_temp[33]_adj_342 (Add_add_temp_adj_2483[33]), .\Add_add_temp[32]_adj_343 (Add_add_temp_adj_2483[32]), 
            .\Add_add_temp[31]_adj_344 (Add_add_temp_adj_2483[31]), .\Add_add_temp[30]_adj_345 (Add_add_temp_adj_2483[30]), 
            .\Add_add_temp[29]_adj_346 (Add_add_temp_adj_2483[29]), .\Add_add_temp[28]_adj_347 (Add_add_temp_adj_2483[28]), 
            .\Add_add_temp[27]_adj_348 (Add_add_temp_adj_2483[27]), .\Add_add_temp[26]_adj_349 (Add_add_temp_adj_2483[26]), 
            .\Add_add_temp[25]_adj_350 (Add_add_temp_adj_2483[25]), .\Add_add_temp[24]_adj_351 (Add_add_temp_adj_2483[24]), 
            .\Add_add_temp[23]_adj_352 (Add_add_temp_adj_2483[23]), .\Add_add_temp[22]_adj_353 (Add_add_temp_adj_2483[22]), 
            .\Add_add_temp[21]_adj_354 (Add_add_temp_adj_2483[21]), .\Add_add_temp[20]_adj_355 (Add_add_temp_adj_2483[20]), 
            .\Add_add_temp[19]_adj_356 (Add_add_temp_adj_2483[19]), .\Add_add_temp[18]_adj_357 (Add_add_temp_adj_2483[18]), 
            .\Add_add_temp[17]_adj_358 (Add_add_temp_adj_2483[17]), .\Add_add_temp[16]_adj_359 (Add_add_temp_adj_2483[16]), 
            .\Add_add_temp[15]_adj_360 (Add_add_temp_adj_2483[15]), .\Add_add_temp[14]_adj_361 (Add_add_temp_adj_2483[14]), 
            .\Add_add_temp[13]_adj_362 (Add_add_temp_adj_2483[13]), .\Add_add_temp[12]_adj_363 (Add_add_temp_adj_2483[12]), 
            .\Add_add_temp[11]_adj_364 (Add_add_temp_adj_2483[11]), .\Add_add_temp[10]_adj_365 (Add_add_temp_adj_2483[10]), 
            .\Add_add_temp[9]_adj_366 (Add_add_temp_adj_2483[9]), .\Add_add_temp[8]_adj_367 (Add_add_temp_adj_2483[8]), 
            .\Add_add_temp[7]_adj_368 (Add_add_temp_adj_2483[7]), .\Add_add_temp[6]_adj_369 (Add_add_temp_adj_2483[6]), 
            .\Add_add_temp[5]_adj_370 (Add_add_temp_adj_2483[5]), .\Add_add_temp[4]_adj_371 (Add_add_temp_adj_2483[4]), 
            .n14328(n14328), .n14327(n14327), .n14326(n14326), .n14322(n14322), 
            .n793_adj_372(n793), .n14325(n14325), .n19782(n19782), .n14324(n14324), 
            .n14323(n14323), .n14321(n14321), .Saturate_out1_31__N_267_adj_373(Saturate_out1_31__N_267), 
            .Saturate_out1_31__N_266_adj_374(Saturate_out1_31__N_266)) /* synthesis lattice_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(55[23] 70[2])
    SB_LUT4 i12403_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[23]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14338));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12403_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12418_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[6]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14353));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12418_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12434_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[22]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14369));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12434_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12435_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[23]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14370));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12435_3_lut.LUT_INIT = 16'haeae;
    SB_IO pin7_pad (.PACKAGE_PIN(pin7), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin7_pad.PIN_TYPE = 6'b101001;
    defparam pin7_pad.PULLUP = 1'b0;
    defparam pin7_pad.NEG_TRIGGER = 1'b0;
    defparam pin7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin8_pad (.PACKAGE_PIN(pin8), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin8_pad.PIN_TYPE = 6'b101001;
    defparam pin8_pad.PULLUP = 1'b0;
    defparam pin8_pad.NEG_TRIGGER = 1'b0;
    defparam pin8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin9_pad (.PACKAGE_PIN(pin9), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin9_pad.PIN_TYPE = 6'b101001;
    defparam pin9_pad.PULLUP = 1'b0;
    defparam pin9_pad.NEG_TRIGGER = 1'b0;
    defparam pin9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i12404_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[24]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14339));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12404_3_lut.LUT_INIT = 16'haeae;
    SB_IO pin10_pad (.PACKAGE_PIN(pin10), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin10_pad.PIN_TYPE = 6'b101001;
    defparam pin10_pad.PULLUP = 1'b0;
    defparam pin10_pad.NEG_TRIGGER = 1'b0;
    defparam pin10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin11_pad (.PACKAGE_PIN(pin11), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin11_pad.PIN_TYPE = 6'b101001;
    defparam pin11_pad.PULLUP = 1'b0;
    defparam pin11_pad.NEG_TRIGGER = 1'b0;
    defparam pin11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin12_pad (.PACKAGE_PIN(pin12), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin12_pad.PIN_TYPE = 6'b101001;
    defparam pin12_pad.PULLUP = 1'b0;
    defparam pin12_pad.NEG_TRIGGER = 1'b0;
    defparam pin12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin13_pad (.PACKAGE_PIN(pin13), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin13_pad.PIN_TYPE = 6'b101001;
    defparam pin13_pad.PULLUP = 1'b0;
    defparam pin13_pad.NEG_TRIGGER = 1'b0;
    defparam pin13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin14_sdo_pad (.PACKAGE_PIN(pin14_sdo), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin14_sdo_pad.PIN_TYPE = 6'b101001;
    defparam pin14_sdo_pad.PULLUP = 1'b0;
    defparam pin14_sdo_pad.NEG_TRIGGER = 1'b0;
    defparam pin14_sdo_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin15_sdi_pad (.PACKAGE_PIN(pin15_sdi), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin15_sdi_pad.PIN_TYPE = 6'b101001;
    defparam pin15_sdi_pad.PULLUP = 1'b0;
    defparam pin15_sdi_pad.NEG_TRIGGER = 1'b0;
    defparam pin15_sdi_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin16_sck_pad (.PACKAGE_PIN(pin16_sck), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin16_sck_pad.PIN_TYPE = 6'b101001;
    defparam pin16_sck_pad.PULLUP = 1'b0;
    defparam pin16_sck_pad.NEG_TRIGGER = 1'b0;
    defparam pin16_sck_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin17_ss_pad (.PACKAGE_PIN(pin17_ss), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin17_ss_pad.PIN_TYPE = 6'b101001;
    defparam pin17_ss_pad.PULLUP = 1'b0;
    defparam pin17_ss_pad.NEG_TRIGGER = 1'b0;
    defparam pin17_ss_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin18_pad (.PACKAGE_PIN(pin18), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin18_pad.PIN_TYPE = 6'b101001;
    defparam pin18_pad.PULLUP = 1'b0;
    defparam pin18_pad.NEG_TRIGGER = 1'b0;
    defparam pin18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin19_pad (.PACKAGE_PIN(pin19), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin19_pad.PIN_TYPE = 6'b101001;
    defparam pin19_pad.PULLUP = 1'b0;
    defparam pin19_pad.NEG_TRIGGER = 1'b0;
    defparam pin19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin20_pad (.PACKAGE_PIN(pin20), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin20_pad.PIN_TYPE = 6'b101001;
    defparam pin20_pad.PULLUP = 1'b0;
    defparam pin20_pad.NEG_TRIGGER = 1'b0;
    defparam pin20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin21_pad (.PACKAGE_PIN(pin21), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin21_pad.PIN_TYPE = 6'b101001;
    defparam pin21_pad.PULLUP = 1'b0;
    defparam pin21_pad.NEG_TRIGGER = 1'b0;
    defparam pin21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin22_pad (.PACKAGE_PIN(pin22), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin22_pad.PIN_TYPE = 6'b101001;
    defparam pin22_pad.PULLUP = 1'b0;
    defparam pin22_pad.NEG_TRIGGER = 1'b0;
    defparam pin22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin23_pad (.PACKAGE_PIN(pin23), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin23_pad.PIN_TYPE = 6'b101001;
    defparam pin23_pad.PULLUP = 1'b0;
    defparam pin23_pad.NEG_TRIGGER = 1'b0;
    defparam pin23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO pin24_pad (.PACKAGE_PIN(pin24), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam pin24_pad.PIN_TYPE = 6'b101001;
    defparam pin24_pad.PULLUP = 1'b0;
    defparam pin24_pad.NEG_TRIGGER = 1'b0;
    defparam pin24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO pin3_clk_16mhz_pad (.PACKAGE_PIN(pin3_clk_16mhz), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(pin3_clk_16mhz_N));   // verilog/TinyFPGA_B.v(4[9:23])
    defparam pin3_clk_16mhz_pad.PIN_TYPE = 6'b000001;
    defparam pin3_clk_16mhz_pad.PULLUP = 1'b0;
    defparam pin3_clk_16mhz_pad.NEG_TRIGGER = 1'b0;
    defparam pin3_clk_16mhz_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i12436_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[24]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14371));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12436_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12405_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[25]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14340));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12405_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12406_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[26]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14341));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12406_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12407_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[27]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14342));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12407_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12437_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[25]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14372));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12437_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12419_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[7]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14354));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12419_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12438_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[26]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14373));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12438_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12408_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[28]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14343));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12408_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12409_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[29]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14344));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12409_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12410_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[30]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14345));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12410_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12439_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[27]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14374));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12439_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12440_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[28]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14375));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12440_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12441_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[29]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14376));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12441_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12411_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[31]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14346));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12411_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12442_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[30]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14377));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12442_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12443_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[31]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14378));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12443_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12444_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[32]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14379));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12444_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12445_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[33]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14380));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12445_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12412_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[32]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14347));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12412_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12413_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[33]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14348));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12413_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12420_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[8]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14355));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12420_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_3_lut (.I0(Saturate_out1_31__N_267_adj_2418), .I1(Saturate_out1_31__N_266_adj_2417), 
            .I2(Add_add_temp_adj_2514[4]), .I3(GND_net), .O(n19765));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12386_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[6]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14321));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12386_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i12414_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[34]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14349));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12414_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i12388_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[8]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14323));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12388_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i11567_4_lut_4_lut (.I0(GND_net), .I1(Look_Up_Table_out1_1[14]), 
            .I2(n628), .I3(Look_Up_Table_out1_1[13]), .O(n4));
    defparam i11567_4_lut_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i12394_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[14]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14329));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12394_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(GND_net), .I1(Look_Up_Table_out1_1[14]), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Amp25_out1[14]), .O(n142));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf888;
    SB_LUT4 i12389_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[9]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14324));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12389_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i1_3_lut_4_lut (.I0(Amp25_out1[14]), .I1(Look_Up_Table_out1_1[15]), 
            .I2(Look_Up_Table_out1_1[14]), .I3(GND_net), .O(n794));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8f88;
    SB_LUT4 i1_3_lut_adj_314 (.I0(Saturate_out1_31__N_267), .I1(Saturate_out1_31__N_266), 
            .I2(Add_add_temp_adj_2483[4]), .I3(GND_net), .O(n19782));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i1_3_lut_adj_314.LUT_INIT = 16'hfefe;
    SB_LUT4 i12390_3_lut (.I0(Saturate_out1_31__N_266), .I1(Add_add_temp_adj_2483[10]), 
            .I2(Saturate_out1_31__N_267), .I3(GND_net), .O(n14325));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12390_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_315 (.I0(GND_net), .I1(Error_sub_temp[30]), .I2(GND_net), 
            .I3(GND_net), .O(n793));
    defparam i1_2_lut_adj_315.LUT_INIT = 16'h2222;
    SB_LUT4 i12680_3_lut (.I0(n146_adj_2423), .I1(Error_sub_temp_adj_2497[30]), 
            .I2(GND_net), .I3(GND_net), .O(n794_adj_2425));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(49[22:38])
    defparam i12680_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i1_2_lut_4_lut (.I0(Amp25_out1[14]), .I1(Error_sub_temp_adj_2497[31]), 
            .I2(GND_net), .I3(Error_sub_temp_adj_2497[30]), .O(n142_adj_2422));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hf888;
    SB_LUT4 i12446_3_lut (.I0(Saturate_out1_31__N_266_adj_2417), .I1(Add_add_temp_adj_2514[34]), 
            .I2(Saturate_out1_31__N_267_adj_2418), .I3(GND_net), .O(n14381));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    defparam i12446_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i1_2_lut_3_lut (.I0(GND_net), .I1(Error_sub_temp[31]), .I2(Error_sub_temp[30]), 
            .I3(GND_net), .O(n142_adj_2419));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he4e4;
    VCC i17141 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module FOC_Current_Control
//

module FOC_Current_Control (Phase_Voltage_0, pin3_clk_16mhz_N_keep, Phase_Voltage_1, 
            Phase_Voltage_2, GND_net, \Amp25_out1[14] , \Product_mul_temp[26] , 
            \Look_Up_Table_out1_1[15] , \Look_Up_Table_out1_1[14] , \Look_Up_Table_out1_1[13] , 
            n628, n142, n139, n794, n4, n14381, \Error_sub_temp[31] , 
            n14380, n14379, n14378, n14377, n14376, n14375, n14374, 
            n14373, n14354, n14372, n14371, n14370, n14369, n14353, 
            n14368, n14367, n14366, n14365, n14364, n14363, n14362, 
            n14361, n14360, n14359, n14352, n14358, n146, n14357, 
            n14356, n793, n141, n794_adj_333, \Add_add_temp[34] , 
            \Add_add_temp[33] , \Add_add_temp[32] , \Add_add_temp[31] , 
            \Add_add_temp[30] , \Add_add_temp[29] , \Add_add_temp[28] , 
            \Add_add_temp[27] , \Add_add_temp[26] , \Add_add_temp[25] , 
            \Add_add_temp[24] , \Add_add_temp[23] , \Add_add_temp[22] , 
            \Add_add_temp[21] , \Add_add_temp[20] , \Add_add_temp[19] , 
            \Add_add_temp[18] , \Add_add_temp[17] , \Add_add_temp[16] , 
            \Add_add_temp[15] , \Add_add_temp[14] , \Add_add_temp[13] , 
            \Add_add_temp[12] , \Add_add_temp[11] , \Add_add_temp[10] , 
            \Add_add_temp[9] , \Add_add_temp[8] , \Add_add_temp[7] , \Add_add_temp[6] , 
            \Add_add_temp[5] , \Add_add_temp[4] , \Error_sub_temp[30] , 
            n19765, n14355, n142_adj_334, Saturate_out1_31__N_267, Saturate_out1_31__N_266, 
            \Error_sub_temp[31]_adj_335 , n146_adj_336, n794_adj_337, 
            n141_adj_338, \Error_sub_temp[30]_adj_339 , n142_adj_340, 
            n14349, n14348, n14347, n14346, n14345, n14344, n14343, 
            n14342, n14341, n14340, n14339, n14338, n14320, n14337, 
            n14336, n14335, n14334, n14333, n14332, n14331, n14330, 
            n14329, \Add_add_temp[34]_adj_341 , \Add_add_temp[33]_adj_342 , 
            \Add_add_temp[32]_adj_343 , \Add_add_temp[31]_adj_344 , \Add_add_temp[30]_adj_345 , 
            \Add_add_temp[29]_adj_346 , \Add_add_temp[28]_adj_347 , \Add_add_temp[27]_adj_348 , 
            \Add_add_temp[26]_adj_349 , \Add_add_temp[25]_adj_350 , \Add_add_temp[24]_adj_351 , 
            \Add_add_temp[23]_adj_352 , \Add_add_temp[22]_adj_353 , \Add_add_temp[21]_adj_354 , 
            \Add_add_temp[20]_adj_355 , \Add_add_temp[19]_adj_356 , \Add_add_temp[18]_adj_357 , 
            \Add_add_temp[17]_adj_358 , \Add_add_temp[16]_adj_359 , \Add_add_temp[15]_adj_360 , 
            \Add_add_temp[14]_adj_361 , \Add_add_temp[13]_adj_362 , \Add_add_temp[12]_adj_363 , 
            \Add_add_temp[11]_adj_364 , \Add_add_temp[10]_adj_365 , \Add_add_temp[9]_adj_366 , 
            \Add_add_temp[8]_adj_367 , \Add_add_temp[7]_adj_368 , \Add_add_temp[6]_adj_369 , 
            \Add_add_temp[5]_adj_370 , \Add_add_temp[4]_adj_371 , n14328, 
            n14327, n14326, n14322, n793_adj_372, n14325, n19782, 
            n14324, n14323, n14321, Saturate_out1_31__N_267_adj_373, 
            Saturate_out1_31__N_266_adj_374) /* synthesis lattice_noprune=1, syn_module_defined=1 */ ;
    output [15:0]Phase_Voltage_0;
    input pin3_clk_16mhz_N_keep;
    output [15:0]Phase_Voltage_1;
    output [15:0]Phase_Voltage_2;
    input GND_net;
    output \Amp25_out1[14] ;
    input \Product_mul_temp[26] ;
    output \Look_Up_Table_out1_1[15] ;
    output \Look_Up_Table_out1_1[14] ;
    output \Look_Up_Table_out1_1[13] ;
    output n628;
    input n142;
    input n139;
    input n794;
    input n4;
    input n14381;
    output \Error_sub_temp[31] ;
    input n14380;
    input n14379;
    input n14378;
    input n14377;
    input n14376;
    input n14375;
    input n14374;
    input n14373;
    input n14354;
    input n14372;
    input n14371;
    input n14370;
    input n14369;
    input n14353;
    input n14368;
    input n14367;
    input n14366;
    input n14365;
    input n14364;
    input n14363;
    input n14362;
    input n14361;
    input n14360;
    input n14359;
    input n14352;
    input n14358;
    output n146;
    input n14357;
    input n14356;
    input n793;
    input n141;
    input n794_adj_333;
    output \Add_add_temp[34] ;
    output \Add_add_temp[33] ;
    output \Add_add_temp[32] ;
    output \Add_add_temp[31] ;
    output \Add_add_temp[30] ;
    output \Add_add_temp[29] ;
    output \Add_add_temp[28] ;
    output \Add_add_temp[27] ;
    output \Add_add_temp[26] ;
    output \Add_add_temp[25] ;
    output \Add_add_temp[24] ;
    output \Add_add_temp[23] ;
    output \Add_add_temp[22] ;
    output \Add_add_temp[21] ;
    output \Add_add_temp[20] ;
    output \Add_add_temp[19] ;
    output \Add_add_temp[18] ;
    output \Add_add_temp[17] ;
    output \Add_add_temp[16] ;
    output \Add_add_temp[15] ;
    output \Add_add_temp[14] ;
    output \Add_add_temp[13] ;
    output \Add_add_temp[12] ;
    output \Add_add_temp[11] ;
    output \Add_add_temp[10] ;
    output \Add_add_temp[9] ;
    output \Add_add_temp[8] ;
    output \Add_add_temp[7] ;
    output \Add_add_temp[6] ;
    output \Add_add_temp[5] ;
    output \Add_add_temp[4] ;
    output \Error_sub_temp[30] ;
    input n19765;
    input n14355;
    input n142_adj_334;
    output Saturate_out1_31__N_267;
    output Saturate_out1_31__N_266;
    output \Error_sub_temp[31]_adj_335 ;
    output n146_adj_336;
    input n794_adj_337;
    input n141_adj_338;
    output \Error_sub_temp[30]_adj_339 ;
    input n142_adj_340;
    input n14349;
    input n14348;
    input n14347;
    input n14346;
    input n14345;
    input n14344;
    input n14343;
    input n14342;
    input n14341;
    input n14340;
    input n14339;
    input n14338;
    input n14320;
    input n14337;
    input n14336;
    input n14335;
    input n14334;
    input n14333;
    input n14332;
    input n14331;
    input n14330;
    input n14329;
    output \Add_add_temp[34]_adj_341 ;
    output \Add_add_temp[33]_adj_342 ;
    output \Add_add_temp[32]_adj_343 ;
    output \Add_add_temp[31]_adj_344 ;
    output \Add_add_temp[30]_adj_345 ;
    output \Add_add_temp[29]_adj_346 ;
    output \Add_add_temp[28]_adj_347 ;
    output \Add_add_temp[27]_adj_348 ;
    output \Add_add_temp[26]_adj_349 ;
    output \Add_add_temp[25]_adj_350 ;
    output \Add_add_temp[24]_adj_351 ;
    output \Add_add_temp[23]_adj_352 ;
    output \Add_add_temp[22]_adj_353 ;
    output \Add_add_temp[21]_adj_354 ;
    output \Add_add_temp[20]_adj_355 ;
    output \Add_add_temp[19]_adj_356 ;
    output \Add_add_temp[18]_adj_357 ;
    output \Add_add_temp[17]_adj_358 ;
    output \Add_add_temp[16]_adj_359 ;
    output \Add_add_temp[15]_adj_360 ;
    output \Add_add_temp[14]_adj_361 ;
    output \Add_add_temp[13]_adj_362 ;
    output \Add_add_temp[12]_adj_363 ;
    output \Add_add_temp[11]_adj_364 ;
    output \Add_add_temp[10]_adj_365 ;
    output \Add_add_temp[9]_adj_366 ;
    output \Add_add_temp[8]_adj_367 ;
    output \Add_add_temp[7]_adj_368 ;
    output \Add_add_temp[6]_adj_369 ;
    output \Add_add_temp[5]_adj_370 ;
    output \Add_add_temp[4]_adj_371 ;
    input n14328;
    input n14327;
    input n14326;
    input n14322;
    input n793_adj_372;
    input n14325;
    input n19782;
    input n14324;
    input n14323;
    input n14321;
    output Saturate_out1_31__N_267_adj_373;
    output Saturate_out1_31__N_266_adj_374;
    
    wire [15:0]svmVoltage_0;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(88[22:34])
    wire [15:0]svmVoltage_1;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(89[22:34])
    wire [15:0]svmVoltage_2;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(90[22:34])
    wire [31:0]abcVoltage_1;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(85[22:34])
    wire [31:0]abcVoltage_2;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(86[22:34])
    wire [15:0]alphaVoltage;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(82[22:34])
    wire [31:0]Gain1_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Clarke_Transform.v(37[22:36])
    wire [15:0]Look_Up_Table_out1_1;   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(77[21:41])
    wire [31:0]dCurrent;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(78[22:30])
    wire [31:0]qCurrent;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(79[22:30])
    wire [15:0]qVoltage;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(81[22:30])
    wire [15:0]dVoltage;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(80[22:30])
    
    wire n610;
    wire [31:0]Product2_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(40[22:39])
    
    wire n86, n576, n414_adj_2204, n267, n218, n236, n120;
    wire [31:0]Product3_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(46[22:39])
    
    wire n26, n71, n138, n44, n89;
    wire [15:0]betaVoltage;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(83[22:33])
    
    wire n209, n19681, n19684, n769, n685, n587, n631, n264, 
        n114, n613, n417, n270, n221, n123, n29, n74, n773, 
        n616, n420_adj_2205, n273, n224, n126, n32, n77, n777, 
        n619, n587_adj_2206, n489, n391, n342, n233, n86_adj_2207, 
        n423, n276, n227, n538, n685_adj_2208, n587_adj_2209, n489_adj_2210, 
        n391_adj_2211, n342_adj_2212, n244, n129, n35, n80, n781, 
        n489_adj_2213, n622, n215, n11, n56, n749, n102, n592, 
        n393, n391_adj_2214, n435, n255, n342_adj_2215, n737, n20, 
        n65, n111, n405, n206, n737_adj_2216, n598, n399, n8, 
        n53, n589, n540, n393_adj_2217, n246, n99, n19351, n50, 
        n741, n592_adj_2218, n543, n396, n249, n102_adj_2219, n8_adj_2220, 
        n53_adj_2221, n745, n595, n546, n399_adj_2222, n252, n105, 
        n11_adj_2223, n56_adj_2224, n749_adj_2225, n598_adj_2226, n549, 
        n402, n255_adj_2227, n108, n14, n59, n753, n601, n552, 
        n405_adj_2228, n258, n111_adj_2229, n17, n62, n757, n604, 
        n555, n408_adj_2230, n261, n114_adj_2231, n20_adj_2232, n65_adj_2233, 
        n761, n607, n558, n411, n264_adj_2234, n117, n23, n68, 
        n765, n610_adj_2235, n561, n414_adj_2236, n267_adj_2237, n761_adj_2238, 
        n120_adj_2239, n26_adj_2240, n71_adj_2241, n769_adj_2242, n613_adj_2243, 
        n564, n417_adj_2244, n17_adj_2245, n62_adj_2246, n601_adj_2247, 
        n244_adj_2248, n288, n195, n239, n408_adj_2249, n108_adj_2250, 
        n402_adj_2251, n270_adj_2252, n745_adj_2253, n141_c, n246_adj_2254, 
        n123_adj_2255, n117_adj_2256, n757_adj_2257, n23_adj_2258, n68_adj_2259, 
        n252_adj_2260, n396_adj_2261, n92, n197, n29_adj_2262, n74_adj_2263, 
        n773_adj_2264, n616_adj_2265, n567, n420_adj_2266, n273_adj_2267, 
        n126_adj_2268, n32_adj_2269, n77_adj_2270, n777_adj_2271, n619_adj_2272, 
        n570, n423_adj_2273, n276_adj_2274, n129_adj_2275, n35_adj_2276, 
        n80_adj_2277, n781_adj_2278, n622_adj_2279, n573, n426_adj_2280, 
        n279, n132, n38, n83, n785, n625, n576_adj_2281, n589_adj_2282, 
        n429, n282, n135, n41, n86_adj_2283, n789, n628_adj_2284, 
        n579, n432_adj_2285, n285, n138_adj_2286, n44_adj_2287, n89_adj_2288, 
        n19604, n685_adj_2289, n587_adj_2290, n631_adj_2291, n538_adj_2292, 
        n582, n489_adj_2293, n391_adj_2294, n435_adj_2295, n342_adj_2296, 
        n244_adj_2297, n288_adj_2298, n195_adj_2299, n141_adj_2300, 
        n92_adj_2301, n203, n99_adj_2302, n19576, n50_adj_2303, n261_adj_2304, 
        n19702, n595_adj_2305, n249_adj_2306, n741_adj_2307, Out_31__N_333;
    wire [31:0]preSatVoltage;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(55[22:35])
    
    wire Out_31__N_332, n426_adj_2308, n258_adj_2309, n19352, Out_31__N_333_adj_2310;
    wire [31:0]preSatVoltage_adj_2383;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(55[22:35])
    
    wire Out_31__N_332_adj_2312, n411_adj_2313, n14_adj_2314, n59_adj_2315, 
        n200, n753_adj_2316, n105_adj_2317, n765_adj_2318, n607_adj_2319, 
        n212, n604_adj_2320, n279_adj_2321, n230, n132_adj_2322, n38_adj_2323, 
        n83_adj_2324, n785_adj_2325, n625_adj_2326, n429_adj_2327, n282_adj_2331, 
        n233_adj_2332, n135_adj_2333, n41_adj_2334, n86_adj_2335, n789_adj_2336, 
        n628_adj_2337, n432_adj_2338, n285_adj_2339;
    
    SB_DFF Delay_Register_out1_2__i48 (.Q(Phase_Voltage_0[15]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[15]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i47 (.Q(Phase_Voltage_0[14]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[14]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i46 (.Q(Phase_Voltage_0[13]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[13]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i45 (.Q(Phase_Voltage_0[12]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[12]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i44 (.Q(Phase_Voltage_0[11]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[11]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i43 (.Q(Phase_Voltage_0[10]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[10]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i42 (.Q(Phase_Voltage_0[9]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[9]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i41 (.Q(Phase_Voltage_0[8]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[8]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i40 (.Q(Phase_Voltage_0[7]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[7]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i39 (.Q(Phase_Voltage_0[6]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[6]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i38 (.Q(Phase_Voltage_0[5]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[5]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i37 (.Q(Phase_Voltage_0[4]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[4]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i36 (.Q(Phase_Voltage_0[3]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[3]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i35 (.Q(Phase_Voltage_0[2]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[2]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i34 (.Q(Phase_Voltage_0[1]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[1]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i33 (.Q(Phase_Voltage_0[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_0[0]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i32 (.Q(Phase_Voltage_1[15]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[15]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i31 (.Q(Phase_Voltage_1[14]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[14]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i30 (.Q(Phase_Voltage_1[13]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[13]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i29 (.Q(Phase_Voltage_1[12]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[12]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i28 (.Q(Phase_Voltage_1[11]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[11]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i27 (.Q(Phase_Voltage_1[10]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[10]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i26 (.Q(Phase_Voltage_1[9]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[9]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i25 (.Q(Phase_Voltage_1[8]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[8]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i24 (.Q(Phase_Voltage_1[7]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[7]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i23 (.Q(Phase_Voltage_1[6]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[6]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i22 (.Q(Phase_Voltage_1[5]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[5]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i1 (.Q(Phase_Voltage_2[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[0]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i21 (.Q(Phase_Voltage_1[4]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[4]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i20 (.Q(Phase_Voltage_1[3]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[3]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i19 (.Q(Phase_Voltage_1[2]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[2]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i18 (.Q(Phase_Voltage_1[1]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[1]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i17 (.Q(Phase_Voltage_1[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_1[0]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i16 (.Q(Phase_Voltage_2[15]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[15]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i15 (.Q(Phase_Voltage_2[14]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[14]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i14 (.Q(Phase_Voltage_2[13]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[13]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i13 (.Q(Phase_Voltage_2[12]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[12]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i12 (.Q(Phase_Voltage_2[11]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[11]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i11 (.Q(Phase_Voltage_2[10]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[10]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i10 (.Q(Phase_Voltage_2[9]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[9]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i9 (.Q(Phase_Voltage_2[8]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[8]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i8 (.Q(Phase_Voltage_2[7]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[7]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i7 (.Q(Phase_Voltage_2[6]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[6]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i6 (.Q(Phase_Voltage_2[5]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[5]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i5 (.Q(Phase_Voltage_2[4]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[4]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i4 (.Q(Phase_Voltage_2[3]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[3]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i3 (.Q(Phase_Voltage_2[2]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[2]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    SB_DFF Delay_Register_out1_2__i2 (.Q(Phase_Voltage_2[1]), .C(pin3_clk_16mhz_N_keep), 
           .D(svmVoltage_2[1]));   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(159[10] 173[8])
    Space_Vector_Modulation u_Space_Vector_Modulation (.svmVoltage_1({svmVoltage_1}), 
            .\abcVoltage_1[31] (abcVoltage_1[31]), .GND_net(GND_net), .\abcVoltage_1[30] (abcVoltage_1[30]), 
            .\abcVoltage_1[29] (abcVoltage_1[29]), .\abcVoltage_1[28] (abcVoltage_1[28]), 
            .\abcVoltage_1[27] (abcVoltage_1[27]), .\abcVoltage_1[26] (abcVoltage_1[26]), 
            .\abcVoltage_1[25] (abcVoltage_1[25]), .\abcVoltage_1[24] (abcVoltage_1[24]), 
            .\abcVoltage_1[23] (abcVoltage_1[23]), .\abcVoltage_1[22] (abcVoltage_1[22]), 
            .\abcVoltage_1[21] (abcVoltage_1[21]), .\abcVoltage_1[20] (abcVoltage_1[20]), 
            .\abcVoltage_1[19] (abcVoltage_1[19]), .\abcVoltage_1[18] (abcVoltage_1[18]), 
            .\abcVoltage_1[17] (abcVoltage_1[17]), .\abcVoltage_1[16] (abcVoltage_1[16]), 
            .svmVoltage_2({svmVoltage_2}), .\abcVoltage_2[31] (abcVoltage_2[31]), 
            .\abcVoltage_2[30] (abcVoltage_2[30]), .\abcVoltage_2[29] (abcVoltage_2[29]), 
            .\abcVoltage_2[28] (abcVoltage_2[28]), .\abcVoltage_2[27] (abcVoltage_2[27]), 
            .\abcVoltage_2[26] (abcVoltage_2[26]), .\abcVoltage_2[25] (abcVoltage_2[25]), 
            .\abcVoltage_2[24] (abcVoltage_2[24]), .\abcVoltage_2[23] (abcVoltage_2[23]), 
            .\abcVoltage_2[22] (abcVoltage_2[22]), .\abcVoltage_2[21] (abcVoltage_2[21]), 
            .\abcVoltage_2[20] (abcVoltage_2[20]), .\abcVoltage_2[19] (abcVoltage_2[19]), 
            .\abcVoltage_2[18] (abcVoltage_2[18]), .\abcVoltage_2[17] (abcVoltage_2[17]), 
            .\abcVoltage_2[16] (abcVoltage_2[16]), .svmVoltage_0({svmVoltage_0}), 
            .alphaVoltage({alphaVoltage}), .\Gain1_mul_temp[2] (Gain1_mul_temp[2]), 
            .\Gain1_mul_temp[1] (Gain1_mul_temp[1]), .\abcVoltage_1[15] (abcVoltage_1[15]), 
            .\abcVoltage_2[15] (abcVoltage_2[15]), .\Gain1_mul_temp[3] (Gain1_mul_temp[3]), 
            .\Gain1_mul_temp[12] (Gain1_mul_temp[12]), .\abcVoltage_2[12] (abcVoltage_2[12]), 
            .\abcVoltage_2[11] (abcVoltage_2[11]), .\abcVoltage_2[8] (abcVoltage_2[8]), 
            .\abcVoltage_2[6] (abcVoltage_2[6]), .\abcVoltage_2[7] (abcVoltage_2[7]), 
            .\abcVoltage_2[3] (abcVoltage_2[3]), .\abcVoltage_2[1] (abcVoltage_2[1]), 
            .\abcVoltage_2[2] (abcVoltage_2[2]), .\abcVoltage_2[10] (abcVoltage_2[10]), 
            .\abcVoltage_2[5] (abcVoltage_2[5]), .\abcVoltage_2[9] (abcVoltage_2[9]), 
            .\abcVoltage_2[4] (abcVoltage_2[4]), .\abcVoltage_2[13] (abcVoltage_2[13]), 
            .\Gain1_mul_temp[5] (Gain1_mul_temp[5]), .\abcVoltage_2[14] (abcVoltage_2[14]), 
            .\Gain1_mul_temp[9] (Gain1_mul_temp[9]), .\Gain1_mul_temp[10] (Gain1_mul_temp[10]), 
            .\Gain1_mul_temp[13] (Gain1_mul_temp[13]), .\Gain1_mul_temp[7] (Gain1_mul_temp[7]), 
            .\Gain1_mul_temp[6] (Gain1_mul_temp[6]), .\Gain1_mul_temp[8] (Gain1_mul_temp[8]), 
            .\abcVoltage_1[14] (abcVoltage_1[14]), .\Gain1_mul_temp[4] (Gain1_mul_temp[4]), 
            .\Gain1_mul_temp[11] (Gain1_mul_temp[11])) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(145[27] 151[55])
    Sine_Cosine u_Sine_Cosine (.GND_net(GND_net), .\Amp25_out1[14] (\Amp25_out1[14] ), 
            .\Product_mul_temp[26] (\Product_mul_temp[26] ), .Look_Up_Table_out1_1({\Look_Up_Table_out1_1[15] , 
            \Look_Up_Table_out1_1[14] , \Look_Up_Table_out1_1[13] , Look_Up_Table_out1_1[12:0]})) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(101[15] 104[31])
    Park_Transform u_Park_Transform (.GND_net(GND_net), .n628(n628), .n142(n142), 
            .\Product_mul_temp[26] (\Product_mul_temp[26] ), .Look_Up_Table_out1_1({\Look_Up_Table_out1_1[15] , 
            \Look_Up_Table_out1_1[14] , \Look_Up_Table_out1_1[13] , Look_Up_Table_out1_1[12:0]}), 
            .\dCurrent[31] (dCurrent[31]), .\dCurrent[30] (dCurrent[30]), 
            .\dCurrent[29] (dCurrent[29]), .\dCurrent[28] (dCurrent[28]), 
            .\dCurrent[27] (dCurrent[27]), .\dCurrent[26] (dCurrent[26]), 
            .\dCurrent[25] (dCurrent[25]), .\dCurrent[24] (dCurrent[24]), 
            .\dCurrent[23] (dCurrent[23]), .\dCurrent[22] (dCurrent[22]), 
            .\dCurrent[21] (dCurrent[21]), .\dCurrent[20] (dCurrent[20]), 
            .\dCurrent[19] (dCurrent[19]), .\dCurrent[18] (dCurrent[18]), 
            .\dCurrent[17] (dCurrent[17]), .\dCurrent[16] (dCurrent[16]), 
            .\dCurrent[15] (dCurrent[15]), .\dCurrent[14] (dCurrent[14]), 
            .\dCurrent[13] (dCurrent[13]), .\dCurrent[12] (dCurrent[12]), 
            .\dCurrent[11] (dCurrent[11]), .\dCurrent[10] (dCurrent[10]), 
            .\dCurrent[9] (dCurrent[9]), .\dCurrent[8] (dCurrent[8]), .\dCurrent[7] (dCurrent[7]), 
            .\dCurrent[6] (dCurrent[6]), .\dCurrent[5] (dCurrent[5]), .\dCurrent[4] (dCurrent[4]), 
            .\qCurrent[3] (qCurrent[3]), .\dCurrent[3] (dCurrent[3]), .n139(n139), 
            .n794(n794), .\qCurrent[31] (qCurrent[31]), .\qCurrent[30] (qCurrent[30]), 
            .\qCurrent[29] (qCurrent[29]), .\qCurrent[28] (qCurrent[28]), 
            .\qCurrent[27] (qCurrent[27]), .\qCurrent[26] (qCurrent[26]), 
            .\qCurrent[25] (qCurrent[25]), .\qCurrent[24] (qCurrent[24]), 
            .\qCurrent[23] (qCurrent[23]), .\qCurrent[22] (qCurrent[22]), 
            .\qCurrent[21] (qCurrent[21]), .\qCurrent[20] (qCurrent[20]), 
            .\qCurrent[19] (qCurrent[19]), .\qCurrent[18] (qCurrent[18]), 
            .\qCurrent[17] (qCurrent[17]), .\qCurrent[16] (qCurrent[16]), 
            .\qCurrent[15] (qCurrent[15]), .\qCurrent[14] (qCurrent[14]), 
            .\qCurrent[13] (qCurrent[13]), .\qCurrent[12] (qCurrent[12]), 
            .\qCurrent[11] (qCurrent[11]), .\qCurrent[10] (qCurrent[10]), 
            .\qCurrent[9] (qCurrent[9]), .\qCurrent[8] (qCurrent[8]), .\qCurrent[7] (qCurrent[7]), 
            .\qCurrent[6] (qCurrent[6]), .\qCurrent[5] (qCurrent[5]), .\qCurrent[4] (qCurrent[4]), 
            .\Amp25_out1[14] (\Amp25_out1[14] ), .n4(n4)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(106[18] 112[37])
    Inverse_Park_Transform u_Inverse_Park_Transform (.\qVoltage[6] (qVoltage[6]), 
            .Look_Up_Table_out1_1({\Look_Up_Table_out1_1[15] , \Look_Up_Table_out1_1[14] , 
            \Look_Up_Table_out1_1[13] , Look_Up_Table_out1_1[12:0]}), .GND_net(GND_net), 
            .\dVoltage[11] (dVoltage[11]), .\qVoltage[7] (qVoltage[7]), 
            .n610(n610), .\Product_mul_temp[26] (\Product_mul_temp[26] ), 
            .\qVoltage[9] (qVoltage[9]), .\Product2_mul_temp[2] (Product2_mul_temp[2]), 
            .n86(n86), .\dVoltage[6] (dVoltage[6]), .\qVoltage[10] (qVoltage[10]), 
            .n576(n576), .n414(n414_adj_2204), .n267(n267), .n218(n218), 
            .\qVoltage[13] (qVoltage[13]), .\qVoltage[14] (qVoltage[14]), 
            .\qVoltage[12] (qVoltage[12]), .n236(n236), .n120(n120), .\qVoltage[3] (qVoltage[3]), 
            .\dVoltage[10] (dVoltage[10]), .\qVoltage[4] (qVoltage[4]), 
            .\Product3_mul_temp[2] (Product3_mul_temp[2]), .n26(n26), .n71(n71), 
            .n138(n138), .n44(n44), .n89(n89), .\betaVoltage[15] (betaVoltage[15]), 
            .n209(n209), .\betaVoltage[14] (betaVoltage[14]), .n19681(n19681), 
            .n19684(n19684), .n769(n769), .n685(n685), .n587(n587), 
            .n631(n631), .\betaVoltage[13] (betaVoltage[13]), .n264(n264), 
            .n114(n114), .n613(n613), .n417(n417), .\betaVoltage[12] (betaVoltage[12]), 
            .\qVoltage[8] (qVoltage[8]), .n270(n270), .n221(n221), .n123(n123), 
            .n29(n29), .n74(n74), .n773(n773), .n616(n616), .n420(n420_adj_2205), 
            .\betaVoltage[11] (betaVoltage[11]), .n273(n273), .n224(n224), 
            .n126(n126), .n32(n32), .n77(n77), .n777(n777), .n619(n619), 
            .n587_adj_203(n587_adj_2206), .n489(n489), .n391(n391), .n342(n342), 
            .\dVoltage[15] (dVoltage[15]), .n233(n233), .n86_adj_204(n86_adj_2207), 
            .n423(n423), .n276(n276), .n227(n227), .n538(n538), .n685_adj_205(n685_adj_2208), 
            .n587_adj_206(n587_adj_2209), .n489_adj_207(n489_adj_2210), 
            .n391_adj_208(n391_adj_2211), .n342_adj_209(n342_adj_2212), 
            .n244(n244), .n129(n129), .n35(n35), .n80(n80), .n781(n781), 
            .n489_adj_210(n489_adj_2213), .n622(n622), .n215(n215), .n11(n11), 
            .n56(n56), .n749(n749), .\qVoltage[15] (qVoltage[15]), .n102(n102), 
            .n592(n592), .n393(n393), .n391_adj_211(n391_adj_2214), .n435(n435), 
            .n255(n255), .n342_adj_212(n342_adj_2215), .n737(n737), .n20(n20), 
            .n65(n65), .n111(n111), .n405(n405), .n206(n206), .n737_adj_213(n737_adj_2216), 
            .n598(n598), .n399(n399), .n8(n8), .n53(n53), .\dVoltage[9] (dVoltage[9]), 
            .n589(n589), .n540(n540), .n393_adj_214(n393_adj_2217), .n246(n246), 
            .n99(n99), .n19351(n19351), .n50(n50), .n741(n741), .n592_adj_215(n592_adj_2218), 
            .n543(n543), .n396(n396), .n249(n249), .n102_adj_216(n102_adj_2219), 
            .n8_adj_217(n8_adj_2220), .n53_adj_218(n53_adj_2221), .n745(n745), 
            .n595(n595), .n546(n546), .n399_adj_219(n399_adj_2222), .n252(n252), 
            .n105(n105), .n11_adj_220(n11_adj_2223), .n56_adj_221(n56_adj_2224), 
            .n749_adj_222(n749_adj_2225), .n598_adj_223(n598_adj_2226), 
            .n549(n549), .n402(n402), .n255_adj_224(n255_adj_2227), .n108(n108), 
            .n14(n14), .n59(n59), .n753(n753), .n601(n601), .n552(n552), 
            .n405_adj_225(n405_adj_2228), .n258(n258), .n111_adj_226(n111_adj_2229), 
            .n17(n17), .n62(n62), .n757(n757), .n604(n604), .n555(n555), 
            .n408(n408_adj_2230), .n261(n261), .n114_adj_227(n114_adj_2231), 
            .n20_adj_228(n20_adj_2232), .n65_adj_229(n65_adj_2233), .n761(n761), 
            .n607(n607), .n558(n558), .n411(n411), .n264_adj_230(n264_adj_2234), 
            .n117(n117), .n23(n23), .n68(n68), .n765(n765), .n610_adj_231(n610_adj_2235), 
            .n561(n561), .n414_adj_232(n414_adj_2236), .n267_adj_233(n267_adj_2237), 
            .n761_adj_234(n761_adj_2238), .n120_adj_235(n120_adj_2239), 
            .n26_adj_236(n26_adj_2240), .n71_adj_237(n71_adj_2241), .n769_adj_238(n769_adj_2242), 
            .n613_adj_239(n613_adj_2243), .n564(n564), .n417_adj_240(n417_adj_2244), 
            .n17_adj_241(n17_adj_2245), .n62_adj_242(n62_adj_2246), .n601_adj_243(n601_adj_2247), 
            .n244_adj_244(n244_adj_2248), .n288(n288), .n195(n195), .n239(n239), 
            .alphaVoltage({alphaVoltage}), .n408_adj_245(n408_adj_2249), 
            .n108_adj_246(n108_adj_2250), .n402_adj_247(n402_adj_2251), 
            .n270_adj_248(n270_adj_2252), .n745_adj_249(n745_adj_2253), 
            .n141(n141_c), .n246_adj_250(n246_adj_2254), .n123_adj_251(n123_adj_2255), 
            .n117_adj_252(n117_adj_2256), .n757_adj_253(n757_adj_2257), 
            .n23_adj_254(n23_adj_2258), .n68_adj_255(n68_adj_2259), .n252_adj_256(n252_adj_2260), 
            .n396_adj_257(n396_adj_2261), .n92(n92), .n197(n197), .n29_adj_258(n29_adj_2262), 
            .n74_adj_259(n74_adj_2263), .n773_adj_260(n773_adj_2264), .n616_adj_261(n616_adj_2265), 
            .n567(n567), .\dVoltage[5] (dVoltage[5]), .n420_adj_262(n420_adj_2266), 
            .n273_adj_263(n273_adj_2267), .n126_adj_264(n126_adj_2268), 
            .n32_adj_265(n32_adj_2269), .n77_adj_266(n77_adj_2270), .n777_adj_267(n777_adj_2271), 
            .n619_adj_268(n619_adj_2272), .n570(n570), .n423_adj_269(n423_adj_2273), 
            .n276_adj_270(n276_adj_2274), .n129_adj_271(n129_adj_2275), 
            .n35_adj_272(n35_adj_2276), .n80_adj_273(n80_adj_2277), .n781_adj_274(n781_adj_2278), 
            .n622_adj_275(n622_adj_2279), .n573(n573), .n426(n426_adj_2280), 
            .n279(n279), .n132(n132), .n38(n38), .n83(n83), .n785(n785), 
            .n625(n625), .n576_adj_276(n576_adj_2281), .n589_adj_277(n589_adj_2282), 
            .n429(n429), .n282(n282), .n135(n135), .n41(n41), .n86_adj_278(n86_adj_2283), 
            .n789(n789), .n628(n628_adj_2284), .n579(n579), .n432(n432_adj_2285), 
            .n285(n285), .n138_adj_279(n138_adj_2286), .n44_adj_280(n44_adj_2287), 
            .n89_adj_281(n89_adj_2288), .n19604(n19604), .n685_adj_282(n685_adj_2289), 
            .n587_adj_283(n587_adj_2290), .n631_adj_284(n631_adj_2291), 
            .n538_adj_285(n538_adj_2292), .n582(n582), .n489_adj_286(n489_adj_2293), 
            .n391_adj_287(n391_adj_2294), .n435_adj_288(n435_adj_2295), 
            .n342_adj_289(n342_adj_2296), .n244_adj_290(n244_adj_2297), 
            .n288_adj_291(n288_adj_2298), .n195_adj_292(n195_adj_2299), 
            .n141_adj_293(n141_adj_2300), .n92_adj_294(n92_adj_2301), .\betaVoltage[10] (betaVoltage[10]), 
            .n203(n203), .n99_adj_295(n99_adj_2302), .\dVoltage[14] (dVoltage[14]), 
            .\dVoltage[7] (dVoltage[7]), .\dVoltage[3] (dVoltage[3]), .\dVoltage[13] (dVoltage[13]), 
            .\betaVoltage[9] (betaVoltage[9]), .n19576(n19576), .n50_adj_296(n50_adj_2303), 
            .\betaVoltage[8] (betaVoltage[8]), .n261_adj_297(n261_adj_2304), 
            .n19702(n19702), .n595_adj_298(n595_adj_2305), .n249_adj_299(n249_adj_2306), 
            .n741_adj_300(n741_adj_2307), .Out_31__N_333(Out_31__N_333), 
            .\preSatVoltage[10] (preSatVoltage[10]), .Out_31__N_332(Out_31__N_332), 
            .\qVoltage[2] (qVoltage[2]), .\qVoltage[5] (qVoltage[5]), .\dVoltage[8] (dVoltage[8]), 
            .n426_adj_301(n426_adj_2308), .n258_adj_302(n258_adj_2309), 
            .\preSatVoltage[13] (preSatVoltage[13]), .\preSatVoltage[12] (preSatVoltage[12]), 
            .\preSatVoltage[19] (preSatVoltage[19]), .\preSatVoltage[22] (preSatVoltage[22]), 
            .\preSatVoltage[23] (preSatVoltage[23]), .n19352(n19352), .Out_31__N_333_adj_303(Out_31__N_333_adj_2310), 
            .\preSatVoltage[10]_adj_304 (preSatVoltage_adj_2383[10]), .Out_31__N_332_adj_305(Out_31__N_332_adj_2312), 
            .\dVoltage[2] (dVoltage[2]), .n411_adj_306(n411_adj_2313), .n14_adj_307(n14_adj_2314), 
            .n59_adj_308(n59_adj_2315), .n200(n200), .n753_adj_309(n753_adj_2316), 
            .n105_adj_310(n105_adj_2317), .n765_adj_311(n765_adj_2318), 
            .n607_adj_312(n607_adj_2319), .n212(n212), .n604_adj_313(n604_adj_2320), 
            .\betaVoltage[7] (betaVoltage[7]), .\betaVoltage[6] (betaVoltage[6]), 
            .n279_adj_314(n279_adj_2321), .n230(n230), .n132_adj_315(n132_adj_2322), 
            .n38_adj_316(n38_adj_2323), .n83_adj_317(n83_adj_2324), .n785_adj_318(n785_adj_2325), 
            .\dVoltage[12] (dVoltage[12]), .\betaVoltage[5] (betaVoltage[5]), 
            .n625_adj_319(n625_adj_2326), .\betaVoltage[4] (betaVoltage[4]), 
            .\betaVoltage[3] (betaVoltage[3]), .\betaVoltage[2] (betaVoltage[2]), 
            .\Gain1_mul_temp[2] (Gain1_mul_temp[2]), .\Gain1_mul_temp[1] (Gain1_mul_temp[1]), 
            .n429_adj_320(n429_adj_2327), .\preSatVoltage[23]_adj_321 (preSatVoltage_adj_2383[23]), 
            .\preSatVoltage[19]_adj_322 (preSatVoltage_adj_2383[19]), .\preSatVoltage[12]_adj_323 (preSatVoltage_adj_2383[12]), 
            .n282_adj_324(n282_adj_2331), .n233_adj_325(n233_adj_2332), 
            .n135_adj_326(n135_adj_2333), .n41_adj_327(n41_adj_2334), .n86_adj_328(n86_adj_2335), 
            .n789_adj_329(n789_adj_2336), .n628_adj_330(n628_adj_2337), 
            .n432_adj_331(n432_adj_2338), .n285_adj_332(n285_adj_2339)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(126[26] 132[53])
    Inverse_Clarke_Transform u_Inverse_Clarke_Transform (.GND_net(GND_net), 
            .\betaVoltage[7] (betaVoltage[7]), .\betaVoltage[12] (betaVoltage[12]), 
            .\betaVoltage[3] (betaVoltage[3]), .\betaVoltage[14] (betaVoltage[14]), 
            .\betaVoltage[15] (betaVoltage[15]), .alphaVoltage({alphaVoltage}), 
            .\betaVoltage[8] (betaVoltage[8]), .\betaVoltage[10] (betaVoltage[10]), 
            .\betaVoltage[5] (betaVoltage[5]), .\betaVoltage[9] (betaVoltage[9]), 
            .\betaVoltage[4] (betaVoltage[4]), .\betaVoltage[13] (betaVoltage[13]), 
            .\betaVoltage[11] (betaVoltage[11]), .\Gain1_mul_temp[1] (Gain1_mul_temp[1]), 
            .\Gain1_mul_temp[13] (Gain1_mul_temp[13]), .\Gain1_mul_temp[12] (Gain1_mul_temp[12]), 
            .\Gain1_mul_temp[11] (Gain1_mul_temp[11]), .\Gain1_mul_temp[10] (Gain1_mul_temp[10]), 
            .\Gain1_mul_temp[9] (Gain1_mul_temp[9]), .\Gain1_mul_temp[8] (Gain1_mul_temp[8]), 
            .\Gain1_mul_temp[7] (Gain1_mul_temp[7]), .\Gain1_mul_temp[6] (Gain1_mul_temp[6]), 
            .\Gain1_mul_temp[5] (Gain1_mul_temp[5]), .\Gain1_mul_temp[4] (Gain1_mul_temp[4]), 
            .\Gain1_mul_temp[3] (Gain1_mul_temp[3]), .\betaVoltage[2] (betaVoltage[2]), 
            .\Gain1_mul_temp[2] (Gain1_mul_temp[2]), .\betaVoltage[6] (betaVoltage[6]), 
            .\abcVoltage_1[31] (abcVoltage_1[31]), .\abcVoltage_1[30] (abcVoltage_1[30]), 
            .\abcVoltage_1[29] (abcVoltage_1[29]), .\abcVoltage_1[28] (abcVoltage_1[28]), 
            .\abcVoltage_1[27] (abcVoltage_1[27]), .\abcVoltage_1[26] (abcVoltage_1[26]), 
            .\abcVoltage_1[25] (abcVoltage_1[25]), .\abcVoltage_1[24] (abcVoltage_1[24]), 
            .\abcVoltage_1[23] (abcVoltage_1[23]), .\abcVoltage_1[22] (abcVoltage_1[22]), 
            .\abcVoltage_1[21] (abcVoltage_1[21]), .\abcVoltage_1[20] (abcVoltage_1[20]), 
            .\abcVoltage_1[19] (abcVoltage_1[19]), .\abcVoltage_1[18] (abcVoltage_1[18]), 
            .\abcVoltage_1[17] (abcVoltage_1[17]), .\abcVoltage_1[16] (abcVoltage_1[16]), 
            .\abcVoltage_1[15] (abcVoltage_1[15]), .\abcVoltage_1[14] (abcVoltage_1[14]), 
            .\abcVoltage_2[31] (abcVoltage_2[31]), .\abcVoltage_2[30] (abcVoltage_2[30]), 
            .\abcVoltage_2[29] (abcVoltage_2[29]), .\abcVoltage_2[28] (abcVoltage_2[28]), 
            .\abcVoltage_2[27] (abcVoltage_2[27]), .\abcVoltage_2[26] (abcVoltage_2[26]), 
            .\abcVoltage_2[25] (abcVoltage_2[25]), .\abcVoltage_2[24] (abcVoltage_2[24]), 
            .\abcVoltage_2[23] (abcVoltage_2[23]), .\abcVoltage_2[22] (abcVoltage_2[22]), 
            .\abcVoltage_2[21] (abcVoltage_2[21]), .\abcVoltage_2[20] (abcVoltage_2[20]), 
            .\abcVoltage_2[19] (abcVoltage_2[19]), .\abcVoltage_2[18] (abcVoltage_2[18]), 
            .\abcVoltage_2[17] (abcVoltage_2[17]), .\abcVoltage_2[16] (abcVoltage_2[16]), 
            .\abcVoltage_2[15] (abcVoltage_2[15]), .\abcVoltage_2[14] (abcVoltage_2[14]), 
            .\abcVoltage_2[13] (abcVoltage_2[13]), .\abcVoltage_2[12] (abcVoltage_2[12]), 
            .\abcVoltage_2[11] (abcVoltage_2[11]), .\abcVoltage_2[10] (abcVoltage_2[10]), 
            .\abcVoltage_2[9] (abcVoltage_2[9]), .\abcVoltage_2[8] (abcVoltage_2[8]), 
            .\abcVoltage_2[7] (abcVoltage_2[7]), .\abcVoltage_2[6] (abcVoltage_2[6]), 
            .\abcVoltage_2[5] (abcVoltage_2[5]), .\abcVoltage_2[4] (abcVoltage_2[4]), 
            .\abcVoltage_2[3] (abcVoltage_2[3]), .\abcVoltage_2[2] (abcVoltage_2[2]), 
            .\abcVoltage_2[1] (abcVoltage_2[1])) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(134[28] 139[57])
    DQ_Current_Control u_DQ_Current_Control (.GND_net(GND_net), .n14381(n14381), 
            .pin3_clk_16mhz_N_keep(pin3_clk_16mhz_N_keep), .\Product_mul_temp[26] (\Product_mul_temp[26] ), 
            .\Error_sub_temp[31] (\Error_sub_temp[31] ), .\preSatVoltage[10] (preSatVoltage[10]), 
            .Out_31__N_333(Out_31__N_333), .Out_31__N_332(Out_31__N_332), 
            .\qVoltage[8] (qVoltage[8]), .\qVoltage[5] (qVoltage[5]), .\qVoltage[2] (qVoltage[2]), 
            .\qVoltage[12] (qVoltage[12]), .n14380(n14380), .\preSatVoltage[23] (preSatVoltage[23]), 
            .\qVoltage[14] (qVoltage[14]), .\qVoltage[9] (qVoltage[9]), 
            .n14379(n14379), .\preSatVoltage[13] (preSatVoltage[13]), .\preSatVoltage[12] (preSatVoltage[12]), 
            .\qVoltage[4] (qVoltage[4]), .\qVoltage[3] (qVoltage[3]), .\qVoltage[15] (qVoltage[15]), 
            .n14378(n14378), .n14377(n14377), .n14376(n14376), .n14375(n14375), 
            .n14374(n14374), .\qVoltage[6] (qVoltage[6]), .n14373(n14373), 
            .\preSatVoltage[22] (preSatVoltage[22]), .\preSatVoltage[19] (preSatVoltage[19]), 
            .\qVoltage[13] (qVoltage[13]), .\qVoltage[10] (qVoltage[10]), 
            .\qVoltage[7] (qVoltage[7]), .n14354(n14354), .n14372(n14372), 
            .n14371(n14371), .n14370(n14370), .n14369(n14369), .n14353(n14353), 
            .n14368(n14368), .n14367(n14367), .n14366(n14366), .n14365(n14365), 
            .n14364(n14364), .n14363(n14363), .n14362(n14362), .n14361(n14361), 
            .n14360(n14360), .n14359(n14359), .n14352(n14352), .n14358(n14358), 
            .\Amp25_out1[14] (\Amp25_out1[14] ), .n146(n146), .n14357(n14357), 
            .n14356(n14356), .n793(n793), .n141(n141), .n794(n794_adj_333), 
            .\Add_add_temp[34] (\Add_add_temp[34] ), .\Add_add_temp[33] (\Add_add_temp[33] ), 
            .\Add_add_temp[32] (\Add_add_temp[32] ), .\Add_add_temp[31] (\Add_add_temp[31] ), 
            .\Add_add_temp[30] (\Add_add_temp[30] ), .\Add_add_temp[29] (\Add_add_temp[29] ), 
            .\Add_add_temp[28] (\Add_add_temp[28] ), .\Add_add_temp[27] (\Add_add_temp[27] ), 
            .\Add_add_temp[26] (\Add_add_temp[26] ), .\Add_add_temp[25] (\Add_add_temp[25] ), 
            .\Add_add_temp[24] (\Add_add_temp[24] ), .\Add_add_temp[23] (\Add_add_temp[23] ), 
            .\Add_add_temp[22] (\Add_add_temp[22] ), .\Add_add_temp[21] (\Add_add_temp[21] ), 
            .\Add_add_temp[20] (\Add_add_temp[20] ), .\Add_add_temp[19] (\Add_add_temp[19] ), 
            .\Add_add_temp[18] (\Add_add_temp[18] ), .\Add_add_temp[17] (\Add_add_temp[17] ), 
            .\Add_add_temp[16] (\Add_add_temp[16] ), .\Add_add_temp[15] (\Add_add_temp[15] ), 
            .\Add_add_temp[14] (\Add_add_temp[14] ), .\Add_add_temp[13] (\Add_add_temp[13] ), 
            .\Add_add_temp[12] (\Add_add_temp[12] ), .\Add_add_temp[11] (\Add_add_temp[11] ), 
            .\Add_add_temp[10] (\Add_add_temp[10] ), .\Add_add_temp[9] (\Add_add_temp[9] ), 
            .\Add_add_temp[8] (\Add_add_temp[8] ), .\Add_add_temp[7] (\Add_add_temp[7] ), 
            .\Add_add_temp[6] (\Add_add_temp[6] ), .\Add_add_temp[5] (\Add_add_temp[5] ), 
            .\Add_add_temp[4] (\Add_add_temp[4] ), .\Error_sub_temp[30] (\Error_sub_temp[30] ), 
            .n19765(n19765), .n14355(n14355), .\qCurrent[3] (qCurrent[3]), 
            .\qCurrent[4] (qCurrent[4]), .\qCurrent[5] (qCurrent[5]), .\qCurrent[6] (qCurrent[6]), 
            .\qCurrent[7] (qCurrent[7]), .\qCurrent[8] (qCurrent[8]), .\qCurrent[9] (qCurrent[9]), 
            .\qCurrent[10] (qCurrent[10]), .\qCurrent[11] (qCurrent[11]), 
            .\qCurrent[12] (qCurrent[12]), .\qCurrent[13] (qCurrent[13]), 
            .\qCurrent[14] (qCurrent[14]), .\qCurrent[15] (qCurrent[15]), 
            .\qCurrent[16] (qCurrent[16]), .\qCurrent[17] (qCurrent[17]), 
            .\qCurrent[18] (qCurrent[18]), .\qCurrent[19] (qCurrent[19]), 
            .\qCurrent[20] (qCurrent[20]), .\qCurrent[21] (qCurrent[21]), 
            .\qCurrent[22] (qCurrent[22]), .\qCurrent[23] (qCurrent[23]), 
            .\qCurrent[24] (qCurrent[24]), .\qCurrent[25] (qCurrent[25]), 
            .\qCurrent[26] (qCurrent[26]), .\qCurrent[27] (qCurrent[27]), 
            .\qCurrent[28] (qCurrent[28]), .\qCurrent[29] (qCurrent[29]), 
            .\qCurrent[30] (qCurrent[30]), .\qCurrent[31] (qCurrent[31]), 
            .n142(n142_adj_334), .Saturate_out1_31__N_267(Saturate_out1_31__N_267), 
            .Saturate_out1_31__N_266(Saturate_out1_31__N_266), .Look_Up_Table_out1_1({\Look_Up_Table_out1_1[15] , 
            \Look_Up_Table_out1_1[14] , \Look_Up_Table_out1_1[13] , Look_Up_Table_out1_1[12:0]}), 
            .n579(n579), .n17(n17), .n267(n267_adj_2237), .n120(n120_adj_2239), 
            .n14(n14), .n414(n414_adj_2236), .n11(n11_adj_2223), .n19604(n19604), 
            .n789(n789), .n785(n785), .n781(n781_adj_2278), .n8(n8_adj_2220), 
            .n777(n777_adj_2271), .n19351(n19351), .n773(n773_adj_2264), 
            .n769(n769_adj_2242), .n765(n765), .n270(n270_adj_2252), .n123(n123_adj_2255), 
            .n761(n761), .n757(n757), .n417(n417_adj_2244), .n753(n753), 
            .n749(n749_adj_2225), .n745(n745), .n741(n741), .n737(n737_adj_2216), 
            .n489(n489), .n489_adj_32(n489_adj_2293), .n342(n342), .n342_adj_33(n342_adj_2296), 
            .n246(n246), .n288(n288_adj_2298), .n285(n285), .n282(n282), 
            .n279(n279), .n276(n276_adj_2274), .n273(n273_adj_2267), .n258(n258), 
            .n255(n255_adj_2227), .n252(n252), .n261(n261), .n249(n249), 
            .n44(n44_adj_2287), .n126(n126_adj_2268), .n420(n420_adj_2266), 
            .n129(n129_adj_2275), .n423(n423_adj_2273), .n41(n41), .n86(n86), 
            .n89(n89_adj_2288), .n86_adj_34(n86_adj_2283), .n83(n83), 
            .n80(n80_adj_2277), .n19702(n19702), .n77(n77_adj_2270), .n74(n74_adj_2263), 
            .n38(n38), .n71(n71_adj_2241), .n68(n68), .n65(n65_adj_2233), 
            .n62(n62), .n59(n59), .n56(n56_adj_2224), .n50(n50), .n53(n53_adj_2221), 
            .n92(n92_adj_2301), .n244(n244_adj_2297), .n35(n35_adj_2276), 
            .n195(n195_adj_2299), .n114(n114_adj_2231), .n108(n108), .n102(n102_adj_2219), 
            .n99(n99), .\Product2_mul_temp[2] (Product2_mul_temp[2]), .n141_adj_35(n141_adj_2300), 
            .n105(n105), .n138(n138_adj_2286), .n135(n135), .n132(n132), 
            .n111(n111_adj_2229), .n32(n32_adj_2269), .n538(n538_adj_2292), 
            .n29(n29_adj_2262), .n426(n426_adj_2280), .n685(n685_adj_2289), 
            .n402(n402), .n429(n429), .n432(n432_adj_2285), .n26(n26_adj_2240), 
            .n391(n391), .n23(n23), .n391_adj_36(n391_adj_2294), .n576(n576), 
            .n576_adj_37(n576_adj_2281), .n573(n573), .n570(n570), .n567(n567), 
            .n564(n564), .n405(n405_adj_2228), .n628(n628_adj_2284), .n625(n625), 
            .n622(n622_adj_2279), .n435(n435_adj_2295), .n619(n619_adj_2272), 
            .n616(n616_adj_2265), .n613(n613_adj_2243), .n610(n610_adj_2235), 
            .n607(n607), .n601(n601), .n561(n561), .n598(n598_adj_2226), 
            .n595(n595), .n592(n592_adj_2218), .n589(n589), .n604(n604), 
            .n631(n631_adj_2291), .n558(n558), .n20(n20_adj_2232), .n264(n264_adj_2234), 
            .n117(n117), .n411(n411), .n587(n587_adj_2206), .n587_adj_38(n587_adj_2290), 
            .n582(n582), .n393(n393_adj_2217), .n408(n408_adj_2230), .n555(n555), 
            .n552(n552), .n549(n549), .n396(n396), .n399(n399_adj_2222), 
            .n546(n546), .n543(n543), .n540(n540), .\Error_sub_temp[31]_adj_39 (\Error_sub_temp[31]_adj_335 ), 
            .n146_adj_40(n146_adj_336), .\preSatVoltage[23]_adj_41 (preSatVoltage_adj_2383[23]), 
            .\preSatVoltage[19]_adj_42 (preSatVoltage_adj_2383[19]), .n794_adj_43(n794_adj_337), 
            .\preSatVoltage[12]_adj_44 (preSatVoltage_adj_2383[12]), .n141_adj_45(n141_adj_338), 
            .\Error_sub_temp[30]_adj_46 (\Error_sub_temp[30]_adj_339 ), .Out_31__N_333_adj_47(Out_31__N_333_adj_2310), 
            .Out_31__N_332_adj_48(Out_31__N_332_adj_2312), .\dVoltage[5] (dVoltage[5]), 
            .\dVoltage[2] (dVoltage[2]), .\dVoltage[8] (dVoltage[8]), .\dVoltage[12] (dVoltage[12]), 
            .\dVoltage[15] (dVoltage[15]), .\dVoltage[13] (dVoltage[13]), 
            .\dVoltage[6] (dVoltage[6]), .\dVoltage[9] (dVoltage[9]), .\dVoltage[11] (dVoltage[11]), 
            .\dVoltage[10] (dVoltage[10]), .\dVoltage[7] (dVoltage[7]), 
            .\dVoltage[3] (dVoltage[3]), .\dVoltage[14] (dVoltage[14]), 
            .\preSatVoltage[10]_adj_49 (preSatVoltage_adj_2383[10]), .n142_adj_50(n142_adj_340), 
            .n14349(n14349), .n14348(n14348), .n14347(n14347), .n14346(n14346), 
            .n14345(n14345), .n14344(n14344), .n14343(n14343), .n14342(n14342), 
            .n14341(n14341), .n14340(n14340), .n14339(n14339), .n14338(n14338), 
            .n14320(n14320), .n14337(n14337), .n14336(n14336), .n14335(n14335), 
            .n14334(n14334), .n14333(n14333), .n14332(n14332), .n14331(n14331), 
            .n14330(n14330), .n14329(n14329), .\Add_add_temp[34]_adj_51 (\Add_add_temp[34]_adj_341 ), 
            .\Add_add_temp[33]_adj_52 (\Add_add_temp[33]_adj_342 ), .\Add_add_temp[32]_adj_53 (\Add_add_temp[32]_adj_343 ), 
            .\Add_add_temp[31]_adj_54 (\Add_add_temp[31]_adj_344 ), .\Add_add_temp[30]_adj_55 (\Add_add_temp[30]_adj_345 ), 
            .\Add_add_temp[29]_adj_56 (\Add_add_temp[29]_adj_346 ), .\Add_add_temp[28]_adj_57 (\Add_add_temp[28]_adj_347 ), 
            .\Add_add_temp[27]_adj_58 (\Add_add_temp[27]_adj_348 ), .\Add_add_temp[26]_adj_59 (\Add_add_temp[26]_adj_349 ), 
            .\Add_add_temp[25]_adj_60 (\Add_add_temp[25]_adj_350 ), .\Add_add_temp[24]_adj_61 (\Add_add_temp[24]_adj_351 ), 
            .\Add_add_temp[23]_adj_62 (\Add_add_temp[23]_adj_352 ), .\Add_add_temp[22]_adj_63 (\Add_add_temp[22]_adj_353 ), 
            .\Add_add_temp[21]_adj_64 (\Add_add_temp[21]_adj_354 ), .\Add_add_temp[20]_adj_65 (\Add_add_temp[20]_adj_355 ), 
            .\Add_add_temp[19]_adj_66 (\Add_add_temp[19]_adj_356 ), .\Add_add_temp[18]_adj_67 (\Add_add_temp[18]_adj_357 ), 
            .\Add_add_temp[17]_adj_68 (\Add_add_temp[17]_adj_358 ), .\Add_add_temp[16]_adj_69 (\Add_add_temp[16]_adj_359 ), 
            .\Add_add_temp[15]_adj_70 (\Add_add_temp[15]_adj_360 ), .\Add_add_temp[14]_adj_71 (\Add_add_temp[14]_adj_361 ), 
            .\Add_add_temp[13]_adj_72 (\Add_add_temp[13]_adj_362 ), .\Add_add_temp[12]_adj_73 (\Add_add_temp[12]_adj_363 ), 
            .\Add_add_temp[11]_adj_74 (\Add_add_temp[11]_adj_364 ), .\Add_add_temp[10]_adj_75 (\Add_add_temp[10]_adj_365 ), 
            .\Add_add_temp[9]_adj_76 (\Add_add_temp[9]_adj_366 ), .\Add_add_temp[8]_adj_77 (\Add_add_temp[8]_adj_367 ), 
            .\Add_add_temp[7]_adj_78 (\Add_add_temp[7]_adj_368 ), .\Add_add_temp[6]_adj_79 (\Add_add_temp[6]_adj_369 ), 
            .\Add_add_temp[5]_adj_80 (\Add_add_temp[5]_adj_370 ), .\Add_add_temp[4]_adj_81 (\Add_add_temp[4]_adj_371 ), 
            .n14328(n14328), .n14327(n14327), .n14326(n14326), .n14322(n14322), 
            .n793_adj_82(n793_adj_372), .n14325(n14325), .n19782(n19782), 
            .n14324(n14324), .n14323(n14323), .n14321(n14321), .Saturate_out1_31__N_267_adj_83(Saturate_out1_31__N_267_adj_373), 
            .Saturate_out1_31__N_266_adj_84(Saturate_out1_31__N_266_adj_374), 
            .\dCurrent[3] (dCurrent[3]), .\dCurrent[4] (dCurrent[4]), .\dCurrent[5] (dCurrent[5]), 
            .\dCurrent[6] (dCurrent[6]), .\dCurrent[7] (dCurrent[7]), .\dCurrent[8] (dCurrent[8]), 
            .\dCurrent[9] (dCurrent[9]), .\dCurrent[10] (dCurrent[10]), 
            .\dCurrent[11] (dCurrent[11]), .\dCurrent[12] (dCurrent[12]), 
            .\dCurrent[13] (dCurrent[13]), .\dCurrent[14] (dCurrent[14]), 
            .\dCurrent[15] (dCurrent[15]), .\dCurrent[16] (dCurrent[16]), 
            .\dCurrent[17] (dCurrent[17]), .\dCurrent[18] (dCurrent[18]), 
            .\dCurrent[19] (dCurrent[19]), .\dCurrent[20] (dCurrent[20]), 
            .\dCurrent[21] (dCurrent[21]), .\dCurrent[22] (dCurrent[22]), 
            .\dCurrent[23] (dCurrent[23]), .\dCurrent[24] (dCurrent[24]), 
            .\dCurrent[25] (dCurrent[25]), .\dCurrent[26] (dCurrent[26]), 
            .\dCurrent[27] (dCurrent[27]), .\dCurrent[28] (dCurrent[28]), 
            .\dCurrent[29] (dCurrent[29]), .\dCurrent[30] (dCurrent[30]), 
            .\dCurrent[31] (dCurrent[31]), .n342_adj_85(n342_adj_2212), 
            .n342_adj_86(n342_adj_2215), .n114_adj_87(n114), .n408_adj_88(n408_adj_2249), 
            .n14_adj_89(n14_adj_2314), .n604_adj_90(n604_adj_2320), .n685_adj_91(n685_adj_2208), 
            .n685_adj_92(n685), .n417_adj_93(n417), .n123_adj_94(n123), 
            .n613_adj_95(n613), .n429_adj_96(n429_adj_2327), .n135_adj_97(n135_adj_2333), 
            .n625_adj_98(n625_adj_2326), .n587_adj_99(n587_adj_2209), .n587_adj_100(n587), 
            .n399_adj_101(n399), .n426_adj_102(n426_adj_2308), .n414_adj_103(n414_adj_2204), 
            .n432_adj_104(n432_adj_2338), .n393_adj_105(n393), .n405_adj_106(n405), 
            .n402_adj_107(n402_adj_2251), .n396_adj_108(n396_adj_2261), 
            .n420_adj_109(n420_adj_2205), .n423_adj_110(n423), .n44_adj_111(n44), 
            .n489_adj_112(n489_adj_2210), .n8_adj_113(n8), .n489_adj_114(n489_adj_2213), 
            .n20_adj_115(n20), .n126_adj_116(n126), .n616_adj_117(n616), 
            .n391_adj_118(n391_adj_2211), .n391_adj_119(n391_adj_2214), 
            .n19576(n19576), .n129_adj_120(n129), .n619_adj_121(n619), 
            .n11_adj_122(n11), .n35_adj_123(n35), .n19352(n19352), .n26_adj_124(n26), 
            .\Product3_mul_temp[2] (Product3_mul_temp[2]), .n120_adj_125(n120), 
            .n111_adj_126(n111), .n102_adj_127(n102), .n99_adj_128(n99_adj_2302), 
            .n108_adj_129(n108_adj_2250), .n138_adj_130(n138), .n132_adj_131(n132_adj_2322), 
            .n105_adj_132(n105_adj_2317), .n610_adj_133(n610), .n595_adj_134(n595_adj_2305), 
            .n23_adj_135(n23_adj_2258), .n622_adj_136(n622), .n41_adj_137(n41_adj_2334), 
            .n601_adj_138(n601_adj_2247), .n592_adj_139(n592), .n598_adj_140(n598), 
            .n589_adj_141(n589_adj_2282), .n628_adj_142(n628_adj_2337), 
            .n32_adj_143(n32), .n538_adj_144(n538), .n29_adj_145(n29), 
            .n17_adj_146(n17_adj_2245), .n71_adj_147(n71), .n83_adj_148(n83_adj_2324), 
            .n59_adj_149(n59_adj_2315), .n50_adj_150(n50_adj_2303), .n92_adj_151(n92), 
            .n68_adj_152(n68_adj_2259), .n62_adj_153(n62_adj_2246), .n53_adj_154(n53), 
            .n65_adj_155(n65), .n38_adj_156(n38_adj_2323), .n56_adj_157(n56), 
            .n80_adj_158(n80), .n244_adj_159(n244), .n233(n233_adj_2332), 
            .n200(n200), .n203(n203), .n86_adj_160(n86_adj_2207), .n77_adj_161(n77), 
            .n197(n197), .n239(n239), .n206(n206), .n86_adj_162(n86_adj_2335), 
            .n215(n215), .n89_adj_163(n89), .n74_adj_164(n74), .n227(n227), 
            .n233_adj_165(n233), .n224(n224), .n221(n221), .n209(n209), 
            .n236(n236), .n230(n230), .n244_adj_166(n244_adj_2248), .n212(n212), 
            .n218(n218), .n279_adj_167(n279_adj_2321), .n270_adj_168(n270), 
            .n267_adj_169(n267), .n255_adj_170(n255), .n285_adj_171(n285_adj_2339), 
            .n264_adj_172(n264), .n258_adj_173(n258_adj_2309), .n249_adj_174(n249_adj_2306), 
            .n246_adj_175(n246_adj_2254), .n273_adj_176(n273), .n282_adj_177(n282_adj_2331), 
            .n261_adj_178(n261_adj_2304), .n19681(n19681), .n288_adj_179(n288), 
            .n276_adj_180(n276), .n252_adj_181(n252_adj_2260), .n789_adj_182(n789_adj_2336), 
            .n785_adj_183(n785_adj_2325), .n765_adj_184(n765_adj_2318), 
            .n753_adj_185(n753_adj_2316), .n741_adj_186(n741_adj_2307), 
            .n757_adj_187(n757_adj_2257), .n745_adj_188(n745_adj_2253), 
            .n761_adj_189(n761_adj_2238), .n195_adj_190(n195), .n737_adj_191(n737), 
            .n749_adj_192(n749), .n781_adj_193(n781), .n777_adj_194(n777), 
            .n773_adj_195(n773), .n769_adj_196(n769), .n19684(n19684), 
            .n435_adj_197(n435), .n141_adj_198(n141_c), .n631_adj_199(n631), 
            .n117_adj_200(n117_adj_2256), .n411_adj_201(n411_adj_2313), 
            .n607_adj_202(n607_adj_2319)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(114[22] 124[45])
    
endmodule
//
// Verilog Description of module Space_Vector_Modulation
//

module Space_Vector_Modulation (svmVoltage_1, \abcVoltage_1[31] , GND_net, 
            \abcVoltage_1[30] , \abcVoltage_1[29] , \abcVoltage_1[28] , 
            \abcVoltage_1[27] , \abcVoltage_1[26] , \abcVoltage_1[25] , 
            \abcVoltage_1[24] , \abcVoltage_1[23] , \abcVoltage_1[22] , 
            \abcVoltage_1[21] , \abcVoltage_1[20] , \abcVoltage_1[19] , 
            \abcVoltage_1[18] , \abcVoltage_1[17] , \abcVoltage_1[16] , 
            svmVoltage_2, \abcVoltage_2[31] , \abcVoltage_2[30] , \abcVoltage_2[29] , 
            \abcVoltage_2[28] , \abcVoltage_2[27] , \abcVoltage_2[26] , 
            \abcVoltage_2[25] , \abcVoltage_2[24] , \abcVoltage_2[23] , 
            \abcVoltage_2[22] , \abcVoltage_2[21] , \abcVoltage_2[20] , 
            \abcVoltage_2[19] , \abcVoltage_2[18] , \abcVoltage_2[17] , 
            \abcVoltage_2[16] , svmVoltage_0, alphaVoltage, \Gain1_mul_temp[2] , 
            \Gain1_mul_temp[1] , \abcVoltage_1[15] , \abcVoltage_2[15] , 
            \Gain1_mul_temp[3] , \Gain1_mul_temp[12] , \abcVoltage_2[12] , 
            \abcVoltage_2[11] , \abcVoltage_2[8] , \abcVoltage_2[6] , 
            \abcVoltage_2[7] , \abcVoltage_2[3] , \abcVoltage_2[1] , \abcVoltage_2[2] , 
            \abcVoltage_2[10] , \abcVoltage_2[5] , \abcVoltage_2[9] , 
            \abcVoltage_2[4] , \abcVoltage_2[13] , \Gain1_mul_temp[5] , 
            \abcVoltage_2[14] , \Gain1_mul_temp[9] , \Gain1_mul_temp[10] , 
            \Gain1_mul_temp[13] , \Gain1_mul_temp[7] , \Gain1_mul_temp[6] , 
            \Gain1_mul_temp[8] , \abcVoltage_1[14] , \Gain1_mul_temp[4] , 
            \Gain1_mul_temp[11] ) /* synthesis syn_module_defined=1 */ ;
    output [15:0]svmVoltage_1;
    input \abcVoltage_1[31] ;
    input GND_net;
    input \abcVoltage_1[30] ;
    input \abcVoltage_1[29] ;
    input \abcVoltage_1[28] ;
    input \abcVoltage_1[27] ;
    input \abcVoltage_1[26] ;
    input \abcVoltage_1[25] ;
    input \abcVoltage_1[24] ;
    input \abcVoltage_1[23] ;
    input \abcVoltage_1[22] ;
    input \abcVoltage_1[21] ;
    input \abcVoltage_1[20] ;
    input \abcVoltage_1[19] ;
    input \abcVoltage_1[18] ;
    input \abcVoltage_1[17] ;
    input \abcVoltage_1[16] ;
    output [15:0]svmVoltage_2;
    input \abcVoltage_2[31] ;
    input \abcVoltage_2[30] ;
    input \abcVoltage_2[29] ;
    input \abcVoltage_2[28] ;
    input \abcVoltage_2[27] ;
    input \abcVoltage_2[26] ;
    input \abcVoltage_2[25] ;
    input \abcVoltage_2[24] ;
    input \abcVoltage_2[23] ;
    input \abcVoltage_2[22] ;
    input \abcVoltage_2[21] ;
    input \abcVoltage_2[20] ;
    input \abcVoltage_2[19] ;
    input \abcVoltage_2[18] ;
    input \abcVoltage_2[17] ;
    input \abcVoltage_2[16] ;
    output [15:0]svmVoltage_0;
    input [15:0]alphaVoltage;
    input \Gain1_mul_temp[2] ;
    input \Gain1_mul_temp[1] ;
    input \abcVoltage_1[15] ;
    input \abcVoltage_2[15] ;
    input \Gain1_mul_temp[3] ;
    input \Gain1_mul_temp[12] ;
    input \abcVoltage_2[12] ;
    input \abcVoltage_2[11] ;
    input \abcVoltage_2[8] ;
    input \abcVoltage_2[6] ;
    input \abcVoltage_2[7] ;
    input \abcVoltage_2[3] ;
    input \abcVoltage_2[1] ;
    input \abcVoltage_2[2] ;
    input \abcVoltage_2[10] ;
    input \abcVoltage_2[5] ;
    input \abcVoltage_2[9] ;
    input \abcVoltage_2[4] ;
    input \abcVoltage_2[13] ;
    input \Gain1_mul_temp[5] ;
    input \abcVoltage_2[14] ;
    input \Gain1_mul_temp[9] ;
    input \Gain1_mul_temp[10] ;
    input \Gain1_mul_temp[13] ;
    input \Gain1_mul_temp[7] ;
    input \Gain1_mul_temp[6] ;
    input \Gain1_mul_temp[8] ;
    input \abcVoltage_1[14] ;
    input \Gain1_mul_temp[4] ;
    input \Gain1_mul_temp[11] ;
    
    wire [16:0]n1;
    
    wire n15654, n15655;
    wire [32:0]Add_add_temp;   // ../../hdlcoderFocCurrentFixptHdl/Space_Vector_Modulation.v(43[22:34])
    wire [31:0]Max_out1;   // ../../hdlcoderFocCurrentFixptHdl/Space_Vector_Modulation.v(38[22:30])
    wire [31:0]Min_out1;   // ../../hdlcoderFocCurrentFixptHdl/Space_Vector_Modulation.v(40[22:30])
    
    wire n15554, n15553, n15552, n15551, n15550, n15549, n15548, 
        n15547, n15546, n15545, n15544, n15543, n15542, n15541, 
        n15540, n15539, n15538, n15537, n15536, n15535, n15534, 
        n15533, n15532, n15531, n15530, n15529, n15528, n15527, 
        n15526, n15525, n15524, n15653, n15652, n15651, n15650, 
        n15649, n15648, n15647, n15646, n15645, n15644, n15643, 
        n15642, n15641, n15640, VCC_net, n15639, n15638, n15637, 
        n15636, n15635, n15634, n15633, n15632, n15631, n15630, 
        n15629, n15628, n15627, n15626, n15625, n15624, n15671, 
        n15670, n15669, n15668, n15667, n15666, n15665, n15664, 
        n15663, n15662, n15661, n15660, n15659, n15658, n15657, 
        n15656;
    
    SB_LUT4 sub_70_add_2_17_lut (.I0(GND_net), .I1(\abcVoltage_1[31] ), 
            .I2(n1[16]), .I3(n15654), .O(svmVoltage_1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_17 (.CI(n15654), .I0(\abcVoltage_1[31] ), .I1(n1[16]), 
            .CO(n15655));
    SB_LUT4 add_6160_33_lut (.I0(GND_net), .I1(Max_out1[31]), .I2(Min_out1[31]), 
            .I3(n15554), .O(Add_add_temp[32])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_32_lut (.I0(GND_net), .I1(Max_out1[31]), .I2(Min_out1[31]), 
            .I3(n15553), .O(Add_add_temp[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_32 (.CI(n15553), .I0(Max_out1[31]), .I1(Min_out1[31]), 
            .CO(n15554));
    SB_LUT4 add_6160_31_lut (.I0(GND_net), .I1(Max_out1[30]), .I2(Min_out1[30]), 
            .I3(n15552), .O(Add_add_temp[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_31 (.CI(n15552), .I0(Max_out1[30]), .I1(Min_out1[30]), 
            .CO(n15553));
    SB_LUT4 add_6160_30_lut (.I0(GND_net), .I1(Max_out1[29]), .I2(Min_out1[29]), 
            .I3(n15551), .O(Add_add_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_30 (.CI(n15551), .I0(Max_out1[29]), .I1(Min_out1[29]), 
            .CO(n15552));
    SB_LUT4 add_6160_29_lut (.I0(GND_net), .I1(Max_out1[28]), .I2(Min_out1[28]), 
            .I3(n15550), .O(Add_add_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_29 (.CI(n15550), .I0(Max_out1[28]), .I1(Min_out1[28]), 
            .CO(n15551));
    SB_LUT4 add_6160_28_lut (.I0(GND_net), .I1(Max_out1[27]), .I2(Min_out1[27]), 
            .I3(n15549), .O(Add_add_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_28 (.CI(n15549), .I0(Max_out1[27]), .I1(Min_out1[27]), 
            .CO(n15550));
    SB_LUT4 add_6160_27_lut (.I0(GND_net), .I1(Max_out1[26]), .I2(Min_out1[26]), 
            .I3(n15548), .O(Add_add_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_27 (.CI(n15548), .I0(Max_out1[26]), .I1(Min_out1[26]), 
            .CO(n15549));
    SB_LUT4 add_6160_26_lut (.I0(GND_net), .I1(Max_out1[25]), .I2(Min_out1[25]), 
            .I3(n15547), .O(Add_add_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_26 (.CI(n15547), .I0(Max_out1[25]), .I1(Min_out1[25]), 
            .CO(n15548));
    SB_LUT4 add_6160_25_lut (.I0(GND_net), .I1(Max_out1[24]), .I2(Min_out1[24]), 
            .I3(n15546), .O(Add_add_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_25 (.CI(n15546), .I0(Max_out1[24]), .I1(Min_out1[24]), 
            .CO(n15547));
    SB_LUT4 add_6160_24_lut (.I0(GND_net), .I1(Max_out1[23]), .I2(Min_out1[23]), 
            .I3(n15545), .O(Add_add_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_24 (.CI(n15545), .I0(Max_out1[23]), .I1(Min_out1[23]), 
            .CO(n15546));
    SB_LUT4 add_6160_23_lut (.I0(GND_net), .I1(Max_out1[22]), .I2(Min_out1[22]), 
            .I3(n15544), .O(Add_add_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_23 (.CI(n15544), .I0(Max_out1[22]), .I1(Min_out1[22]), 
            .CO(n15545));
    SB_LUT4 add_6160_22_lut (.I0(GND_net), .I1(Max_out1[21]), .I2(Min_out1[21]), 
            .I3(n15543), .O(Add_add_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_22 (.CI(n15543), .I0(Max_out1[21]), .I1(Min_out1[21]), 
            .CO(n15544));
    SB_LUT4 add_6160_21_lut (.I0(GND_net), .I1(Max_out1[20]), .I2(Min_out1[20]), 
            .I3(n15542), .O(Add_add_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_21 (.CI(n15542), .I0(Max_out1[20]), .I1(Min_out1[20]), 
            .CO(n15543));
    SB_LUT4 add_6160_20_lut (.I0(GND_net), .I1(Max_out1[19]), .I2(Min_out1[19]), 
            .I3(n15541), .O(Add_add_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_20 (.CI(n15541), .I0(Max_out1[19]), .I1(Min_out1[19]), 
            .CO(n15542));
    SB_LUT4 add_6160_19_lut (.I0(GND_net), .I1(Max_out1[18]), .I2(Min_out1[18]), 
            .I3(n15540), .O(Add_add_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_19 (.CI(n15540), .I0(Max_out1[18]), .I1(Min_out1[18]), 
            .CO(n15541));
    SB_LUT4 add_6160_18_lut (.I0(GND_net), .I1(Max_out1[17]), .I2(Min_out1[17]), 
            .I3(n15539), .O(Add_add_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_18 (.CI(n15539), .I0(Max_out1[17]), .I1(Min_out1[17]), 
            .CO(n15540));
    SB_CARRY add_6160_17 (.CI(n15538), .I0(Max_out1[16]), .I1(Min_out1[16]), 
            .CO(n15539));
    SB_CARRY add_6160_16 (.CI(n15537), .I0(Max_out1[15]), .I1(Min_out1[15]), 
            .CO(n15538));
    SB_CARRY add_6160_15 (.CI(n15536), .I0(Max_out1[14]), .I1(Min_out1[14]), 
            .CO(n15537));
    SB_CARRY add_6160_14 (.CI(n15535), .I0(Max_out1[13]), .I1(Min_out1[13]), 
            .CO(n15536));
    SB_CARRY add_6160_13 (.CI(n15534), .I0(Max_out1[12]), .I1(Min_out1[12]), 
            .CO(n15535));
    SB_CARRY add_6160_12 (.CI(n15533), .I0(Max_out1[11]), .I1(Min_out1[11]), 
            .CO(n15534));
    SB_CARRY add_6160_11 (.CI(n15532), .I0(Max_out1[10]), .I1(Min_out1[10]), 
            .CO(n15533));
    SB_CARRY add_6160_10 (.CI(n15531), .I0(Max_out1[9]), .I1(Min_out1[9]), 
            .CO(n15532));
    SB_CARRY add_6160_9 (.CI(n15530), .I0(Max_out1[8]), .I1(Min_out1[8]), 
            .CO(n15531));
    SB_CARRY add_6160_8 (.CI(n15529), .I0(Max_out1[7]), .I1(Min_out1[7]), 
            .CO(n15530));
    SB_CARRY add_6160_7 (.CI(n15528), .I0(Max_out1[6]), .I1(Min_out1[6]), 
            .CO(n15529));
    SB_CARRY add_6160_6 (.CI(n15527), .I0(Max_out1[5]), .I1(Min_out1[5]), 
            .CO(n15528));
    SB_CARRY add_6160_5 (.CI(n15526), .I0(Max_out1[4]), .I1(Min_out1[4]), 
            .CO(n15527));
    SB_CARRY add_6160_4 (.CI(n15525), .I0(Max_out1[3]), .I1(Min_out1[3]), 
            .CO(n15526));
    SB_CARRY add_6160_3 (.CI(n15524), .I0(Max_out1[2]), .I1(Min_out1[2]), 
            .CO(n15525));
    SB_CARRY add_6160_2 (.CI(GND_net), .I0(Max_out1[1]), .I1(Min_out1[1]), 
            .CO(n15524));
    SB_LUT4 sub_69_inv_0_i15_1_lut (.I0(Add_add_temp[31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));
    defparam sub_69_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_70_add_2_16_lut (.I0(GND_net), .I1(\abcVoltage_1[30] ), 
            .I2(n1[14]), .I3(n15653), .O(svmVoltage_1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_16 (.CI(n15653), .I0(\abcVoltage_1[30] ), .I1(n1[14]), 
            .CO(n15654));
    SB_LUT4 sub_70_add_2_15_lut (.I0(GND_net), .I1(\abcVoltage_1[29] ), 
            .I2(n1[13]), .I3(n15652), .O(svmVoltage_1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_15 (.CI(n15652), .I0(\abcVoltage_1[29] ), .I1(n1[13]), 
            .CO(n15653));
    SB_LUT4 sub_70_add_2_14_lut (.I0(GND_net), .I1(\abcVoltage_1[28] ), 
            .I2(n1[12]), .I3(n15651), .O(svmVoltage_1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_14 (.CI(n15651), .I0(\abcVoltage_1[28] ), .I1(n1[12]), 
            .CO(n15652));
    SB_LUT4 sub_70_add_2_13_lut (.I0(GND_net), .I1(\abcVoltage_1[27] ), 
            .I2(n1[11]), .I3(n15650), .O(svmVoltage_1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_13 (.CI(n15650), .I0(\abcVoltage_1[27] ), .I1(n1[11]), 
            .CO(n15651));
    SB_LUT4 sub_70_add_2_12_lut (.I0(GND_net), .I1(\abcVoltage_1[26] ), 
            .I2(n1[10]), .I3(n15649), .O(svmVoltage_1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_12 (.CI(n15649), .I0(\abcVoltage_1[26] ), .I1(n1[10]), 
            .CO(n15650));
    SB_LUT4 sub_70_add_2_11_lut (.I0(GND_net), .I1(\abcVoltage_1[25] ), 
            .I2(n1[9]), .I3(n15648), .O(svmVoltage_1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_11 (.CI(n15648), .I0(\abcVoltage_1[25] ), .I1(n1[9]), 
            .CO(n15649));
    SB_LUT4 sub_70_add_2_10_lut (.I0(GND_net), .I1(\abcVoltage_1[24] ), 
            .I2(n1[8]), .I3(n15647), .O(svmVoltage_1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_10 (.CI(n15647), .I0(\abcVoltage_1[24] ), .I1(n1[8]), 
            .CO(n15648));
    SB_LUT4 sub_70_add_2_9_lut (.I0(GND_net), .I1(\abcVoltage_1[23] ), .I2(n1[7]), 
            .I3(n15646), .O(svmVoltage_1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_9 (.CI(n15646), .I0(\abcVoltage_1[23] ), .I1(n1[7]), 
            .CO(n15647));
    SB_LUT4 sub_70_add_2_8_lut (.I0(GND_net), .I1(\abcVoltage_1[22] ), .I2(n1[6]), 
            .I3(n15645), .O(svmVoltage_1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_8 (.CI(n15645), .I0(\abcVoltage_1[22] ), .I1(n1[6]), 
            .CO(n15646));
    SB_LUT4 sub_70_add_2_7_lut (.I0(GND_net), .I1(\abcVoltage_1[21] ), .I2(n1[5]), 
            .I3(n15644), .O(svmVoltage_1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_7 (.CI(n15644), .I0(\abcVoltage_1[21] ), .I1(n1[5]), 
            .CO(n15645));
    SB_LUT4 sub_70_add_2_6_lut (.I0(GND_net), .I1(\abcVoltage_1[20] ), .I2(n1[4]), 
            .I3(n15643), .O(svmVoltage_1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_6 (.CI(n15643), .I0(\abcVoltage_1[20] ), .I1(n1[4]), 
            .CO(n15644));
    SB_LUT4 sub_70_add_2_5_lut (.I0(GND_net), .I1(\abcVoltage_1[19] ), .I2(n1[3]), 
            .I3(n15642), .O(svmVoltage_1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_5 (.CI(n15642), .I0(\abcVoltage_1[19] ), .I1(n1[3]), 
            .CO(n15643));
    SB_LUT4 sub_70_add_2_4_lut (.I0(GND_net), .I1(\abcVoltage_1[18] ), .I2(n1[2]), 
            .I3(n15641), .O(svmVoltage_1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_4 (.CI(n15641), .I0(\abcVoltage_1[18] ), .I1(n1[2]), 
            .CO(n15642));
    SB_LUT4 sub_70_add_2_3_lut (.I0(GND_net), .I1(\abcVoltage_1[17] ), .I2(n1[1]), 
            .I3(n15640), .O(svmVoltage_1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_70_add_2_3 (.CI(n15640), .I0(\abcVoltage_1[17] ), .I1(n1[1]), 
            .CO(n15641));
    SB_CARRY sub_70_add_2_2 (.CI(VCC_net), .I0(\abcVoltage_1[16] ), .I1(n1[0]), 
            .CO(n15640));
    SB_LUT4 sub_71_add_2_18_lut (.I0(GND_net), .I1(\abcVoltage_2[31] ), 
            .I2(n1[16]), .I3(n15639), .O(svmVoltage_2[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_71_add_2_17_lut (.I0(GND_net), .I1(\abcVoltage_2[31] ), 
            .I2(n1[16]), .I3(n15638), .O(svmVoltage_2[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_17 (.CI(n15638), .I0(\abcVoltage_2[31] ), .I1(n1[16]), 
            .CO(n15639));
    SB_LUT4 sub_69_inv_0_i17_1_lut (.I0(Add_add_temp[32]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));
    defparam sub_69_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_71_add_2_16_lut (.I0(GND_net), .I1(\abcVoltage_2[30] ), 
            .I2(n1[14]), .I3(n15637), .O(svmVoltage_2[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_16 (.CI(n15637), .I0(\abcVoltage_2[30] ), .I1(n1[14]), 
            .CO(n15638));
    SB_LUT4 sub_71_add_2_15_lut (.I0(GND_net), .I1(\abcVoltage_2[29] ), 
            .I2(n1[13]), .I3(n15636), .O(svmVoltage_2[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_15 (.CI(n15636), .I0(\abcVoltage_2[29] ), .I1(n1[13]), 
            .CO(n15637));
    SB_LUT4 sub_71_add_2_14_lut (.I0(GND_net), .I1(\abcVoltage_2[28] ), 
            .I2(n1[12]), .I3(n15635), .O(svmVoltage_2[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_14 (.CI(n15635), .I0(\abcVoltage_2[28] ), .I1(n1[12]), 
            .CO(n15636));
    SB_LUT4 sub_71_add_2_13_lut (.I0(GND_net), .I1(\abcVoltage_2[27] ), 
            .I2(n1[11]), .I3(n15634), .O(svmVoltage_2[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_13 (.CI(n15634), .I0(\abcVoltage_2[27] ), .I1(n1[11]), 
            .CO(n15635));
    SB_LUT4 sub_71_add_2_12_lut (.I0(GND_net), .I1(\abcVoltage_2[26] ), 
            .I2(n1[10]), .I3(n15633), .O(svmVoltage_2[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_12 (.CI(n15633), .I0(\abcVoltage_2[26] ), .I1(n1[10]), 
            .CO(n15634));
    SB_LUT4 sub_71_add_2_11_lut (.I0(GND_net), .I1(\abcVoltage_2[25] ), 
            .I2(n1[9]), .I3(n15632), .O(svmVoltage_2[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_11 (.CI(n15632), .I0(\abcVoltage_2[25] ), .I1(n1[9]), 
            .CO(n15633));
    SB_LUT4 sub_71_add_2_10_lut (.I0(GND_net), .I1(\abcVoltage_2[24] ), 
            .I2(n1[8]), .I3(n15631), .O(svmVoltage_2[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_10 (.CI(n15631), .I0(\abcVoltage_2[24] ), .I1(n1[8]), 
            .CO(n15632));
    SB_LUT4 sub_71_add_2_9_lut (.I0(GND_net), .I1(\abcVoltage_2[23] ), .I2(n1[7]), 
            .I3(n15630), .O(svmVoltage_2[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_9 (.CI(n15630), .I0(\abcVoltage_2[23] ), .I1(n1[7]), 
            .CO(n15631));
    SB_LUT4 sub_71_add_2_8_lut (.I0(GND_net), .I1(\abcVoltage_2[22] ), .I2(n1[6]), 
            .I3(n15629), .O(svmVoltage_2[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_8 (.CI(n15629), .I0(\abcVoltage_2[22] ), .I1(n1[6]), 
            .CO(n15630));
    SB_LUT4 sub_71_add_2_7_lut (.I0(GND_net), .I1(\abcVoltage_2[21] ), .I2(n1[5]), 
            .I3(n15628), .O(svmVoltage_2[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_7 (.CI(n15628), .I0(\abcVoltage_2[21] ), .I1(n1[5]), 
            .CO(n15629));
    SB_LUT4 sub_71_add_2_6_lut (.I0(GND_net), .I1(\abcVoltage_2[20] ), .I2(n1[4]), 
            .I3(n15627), .O(svmVoltage_2[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_6 (.CI(n15627), .I0(\abcVoltage_2[20] ), .I1(n1[4]), 
            .CO(n15628));
    SB_LUT4 sub_71_add_2_5_lut (.I0(GND_net), .I1(\abcVoltage_2[19] ), .I2(n1[3]), 
            .I3(n15626), .O(svmVoltage_2[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_5 (.CI(n15626), .I0(\abcVoltage_2[19] ), .I1(n1[3]), 
            .CO(n15627));
    SB_LUT4 sub_71_add_2_4_lut (.I0(GND_net), .I1(\abcVoltage_2[18] ), .I2(n1[2]), 
            .I3(n15625), .O(svmVoltage_2[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_4 (.CI(n15625), .I0(\abcVoltage_2[18] ), .I1(n1[2]), 
            .CO(n15626));
    SB_LUT4 sub_71_add_2_3_lut (.I0(GND_net), .I1(\abcVoltage_2[17] ), .I2(n1[1]), 
            .I3(n15624), .O(svmVoltage_2[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_71_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_71_add_2_3 (.CI(n15624), .I0(\abcVoltage_2[17] ), .I1(n1[1]), 
            .CO(n15625));
    SB_CARRY sub_71_add_2_2 (.CI(VCC_net), .I0(\abcVoltage_2[16] ), .I1(n1[0]), 
            .CO(n15624));
    SB_LUT4 sub_69_add_2_18_lut (.I0(GND_net), .I1(alphaVoltage[15]), .I2(n1[16]), 
            .I3(n15671), .O(svmVoltage_0[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_17_lut (.I0(GND_net), .I1(alphaVoltage[15]), .I2(n1[16]), 
            .I3(n15670), .O(svmVoltage_0[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_17 (.CI(n15670), .I0(alphaVoltage[15]), .I1(n1[16]), 
            .CO(n15671));
    SB_LUT4 sub_69_add_2_16_lut (.I0(GND_net), .I1(alphaVoltage[15]), .I2(n1[14]), 
            .I3(n15669), .O(svmVoltage_0[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_16 (.CI(n15669), .I0(alphaVoltage[15]), .I1(n1[14]), 
            .CO(n15670));
    SB_LUT4 sub_69_add_2_15_lut (.I0(GND_net), .I1(alphaVoltage[14]), .I2(n1[13]), 
            .I3(n15668), .O(svmVoltage_0[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_15 (.CI(n15668), .I0(alphaVoltage[14]), .I1(n1[13]), 
            .CO(n15669));
    SB_LUT4 sub_69_add_2_14_lut (.I0(GND_net), .I1(alphaVoltage[13]), .I2(n1[12]), 
            .I3(n15667), .O(svmVoltage_0[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_14 (.CI(n15667), .I0(alphaVoltage[13]), .I1(n1[12]), 
            .CO(n15668));
    SB_LUT4 sub_69_add_2_13_lut (.I0(GND_net), .I1(alphaVoltage[12]), .I2(n1[11]), 
            .I3(n15666), .O(svmVoltage_0[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_13 (.CI(n15666), .I0(alphaVoltage[12]), .I1(n1[11]), 
            .CO(n15667));
    SB_LUT4 sub_69_add_2_12_lut (.I0(GND_net), .I1(alphaVoltage[11]), .I2(n1[10]), 
            .I3(n15665), .O(svmVoltage_0[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_12 (.CI(n15665), .I0(alphaVoltage[11]), .I1(n1[10]), 
            .CO(n15666));
    SB_LUT4 sub_69_add_2_11_lut (.I0(GND_net), .I1(alphaVoltage[10]), .I2(n1[9]), 
            .I3(n15664), .O(svmVoltage_0[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_11 (.CI(n15664), .I0(alphaVoltage[10]), .I1(n1[9]), 
            .CO(n15665));
    SB_LUT4 sub_69_add_2_10_lut (.I0(GND_net), .I1(alphaVoltage[9]), .I2(n1[8]), 
            .I3(n15663), .O(svmVoltage_0[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_10 (.CI(n15663), .I0(alphaVoltage[9]), .I1(n1[8]), 
            .CO(n15664));
    SB_LUT4 sub_69_add_2_9_lut (.I0(GND_net), .I1(alphaVoltage[8]), .I2(n1[7]), 
            .I3(n15662), .O(svmVoltage_0[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_9 (.CI(n15662), .I0(alphaVoltage[8]), .I1(n1[7]), 
            .CO(n15663));
    SB_LUT4 sub_69_add_2_8_lut (.I0(GND_net), .I1(alphaVoltage[7]), .I2(n1[6]), 
            .I3(n15661), .O(svmVoltage_0[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_8 (.CI(n15661), .I0(alphaVoltage[7]), .I1(n1[6]), 
            .CO(n15662));
    SB_LUT4 sub_69_add_2_7_lut (.I0(GND_net), .I1(alphaVoltage[6]), .I2(n1[5]), 
            .I3(n15660), .O(svmVoltage_0[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_7 (.CI(n15660), .I0(alphaVoltage[6]), .I1(n1[5]), 
            .CO(n15661));
    SB_LUT4 sub_69_add_2_6_lut (.I0(GND_net), .I1(alphaVoltage[5]), .I2(n1[4]), 
            .I3(n15659), .O(svmVoltage_0[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_6 (.CI(n15659), .I0(alphaVoltage[5]), .I1(n1[4]), 
            .CO(n15660));
    SB_LUT4 sub_69_add_2_5_lut (.I0(GND_net), .I1(alphaVoltage[4]), .I2(n1[3]), 
            .I3(n15658), .O(svmVoltage_0[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_5 (.CI(n15658), .I0(alphaVoltage[4]), .I1(n1[3]), 
            .CO(n15659));
    SB_LUT4 sub_69_add_2_4_lut (.I0(GND_net), .I1(alphaVoltage[3]), .I2(n1[2]), 
            .I3(n15657), .O(svmVoltage_0[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_4 (.CI(n15657), .I0(alphaVoltage[3]), .I1(n1[2]), 
            .CO(n15658));
    SB_LUT4 sub_69_add_2_3_lut (.I0(GND_net), .I1(alphaVoltage[2]), .I2(n1[1]), 
            .I3(n15656), .O(svmVoltage_0[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_3 (.CI(n15656), .I0(alphaVoltage[2]), .I1(n1[1]), 
            .CO(n15657));
    SB_CARRY sub_69_add_2_2 (.CI(VCC_net), .I0(alphaVoltage[1]), .I1(n1[0]), 
            .CO(n15656));
    SB_LUT4 sub_70_add_2_18_lut (.I0(GND_net), .I1(\abcVoltage_1[31] ), 
            .I2(n1[16]), .I3(n15655), .O(svmVoltage_1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_70_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_inv_0_i1_1_lut (.I0(Add_add_temp[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));
    defparam sub_69_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i2_1_lut (.I0(Add_add_temp[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));
    defparam sub_69_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i3_1_lut (.I0(Add_add_temp[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));
    defparam sub_69_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i4_1_lut (.I0(Add_add_temp[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));
    defparam sub_69_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i5_1_lut (.I0(Add_add_temp[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));
    defparam sub_69_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i6_1_lut (.I0(Add_add_temp[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));
    defparam sub_69_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i7_1_lut (.I0(Add_add_temp[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));
    defparam sub_69_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i8_1_lut (.I0(Add_add_temp[24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));
    defparam sub_69_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i9_1_lut (.I0(Add_add_temp[25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));
    defparam sub_69_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i10_1_lut (.I0(Add_add_temp[26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));
    defparam sub_69_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i11_1_lut (.I0(Add_add_temp[27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));
    defparam sub_69_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i12_1_lut (.I0(Add_add_temp[28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));
    defparam sub_69_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i13_1_lut (.I0(Add_add_temp[29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));
    defparam sub_69_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_69_inv_0_i14_1_lut (.I0(Add_add_temp[30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));
    defparam sub_69_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    Min u_Min (.\abcVoltage_1[30] (\abcVoltage_1[30] ), .alphaVoltage({alphaVoltage}), 
        .GND_net(GND_net), .\Gain1_mul_temp[2] (\Gain1_mul_temp[2] ), .\Gain1_mul_temp[1] (\Gain1_mul_temp[1] ), 
        .\abcVoltage_1[26] (\abcVoltage_1[26] ), .\abcVoltage_2[26] (\abcVoltage_2[26] ), 
        .\abcVoltage_1[29] (\abcVoltage_1[29] ), .\abcVoltage_2[29] (\abcVoltage_2[29] ), 
        .\abcVoltage_1[28] (\abcVoltage_1[28] ), .\abcVoltage_2[28] (\abcVoltage_2[28] ), 
        .\abcVoltage_1[27] (\abcVoltage_1[27] ), .\abcVoltage_2[27] (\abcVoltage_2[27] ), 
        .\abcVoltage_1[19] (\abcVoltage_1[19] ), .\abcVoltage_2[19] (\abcVoltage_2[19] ), 
        .\abcVoltage_1[21] (\abcVoltage_1[21] ), .\abcVoltage_1[20] (\abcVoltage_1[20] ), 
        .\abcVoltage_2[20] (\abcVoltage_2[20] ), .\abcVoltage_2[21] (\abcVoltage_2[21] ), 
        .\abcVoltage_1[16] (\abcVoltage_1[16] ), .\abcVoltage_1[15] (\abcVoltage_1[15] ), 
        .\abcVoltage_2[15] (\abcVoltage_2[15] ), .\abcVoltage_2[16] (\abcVoltage_2[16] ), 
        .\Gain1_mul_temp[3] (\Gain1_mul_temp[3] ), .\abcVoltage_1[18] (\abcVoltage_1[18] ), 
        .\abcVoltage_2[18] (\abcVoltage_2[18] ), .\abcVoltage_1[17] (\abcVoltage_1[17] ), 
        .\abcVoltage_2[17] (\abcVoltage_2[17] ), .\abcVoltage_1[25] (\abcVoltage_1[25] ), 
        .\abcVoltage_1[23] (\abcVoltage_1[23] ), .\abcVoltage_1[24] (\abcVoltage_1[24] ), 
        .\abcVoltage_2[23] (\abcVoltage_2[23] ), .\abcVoltage_2[24] (\abcVoltage_2[24] ), 
        .\abcVoltage_2[25] (\abcVoltage_2[25] ), .\abcVoltage_1[22] (\abcVoltage_1[22] ), 
        .\Gain1_mul_temp[12] (\Gain1_mul_temp[12] ), .\abcVoltage_2[12] (\abcVoltage_2[12] ), 
        .\abcVoltage_2[22] (\abcVoltage_2[22] ), .\abcVoltage_1[31] (\abcVoltage_1[31] ), 
        .\abcVoltage_2[11] (\abcVoltage_2[11] ), .\abcVoltage_2[8] (\abcVoltage_2[8] ), 
        .\abcVoltage_2[6] (\abcVoltage_2[6] ), .\abcVoltage_2[7] (\abcVoltage_2[7] ), 
        .\abcVoltage_2[3] (\abcVoltage_2[3] ), .\abcVoltage_2[1] (\abcVoltage_2[1] ), 
        .\Min_out1[1] (Min_out1[1]), .\abcVoltage_2[2] (\abcVoltage_2[2] ), 
        .\Min_out1[2] (Min_out1[2]), .\Min_out1[3] (Min_out1[3]), .\abcVoltage_2[10] (\abcVoltage_2[10] ), 
        .\abcVoltage_2[5] (\abcVoltage_2[5] ), .\abcVoltage_2[9] (\abcVoltage_2[9] ), 
        .\abcVoltage_2[4] (\abcVoltage_2[4] ), .\abcVoltage_2[13] (\abcVoltage_2[13] ), 
        .\Gain1_mul_temp[5] (\Gain1_mul_temp[5] ), .\abcVoltage_2[14] (\abcVoltage_2[14] ), 
        .\Min_out1[5] (Min_out1[5]), .\Min_out1[15] (Min_out1[15]), .\Min_out1[16] (Min_out1[16]), 
        .\Min_out1[17] (Min_out1[17]), .\Min_out1[18] (Min_out1[18]), .\abcVoltage_2[30] (\abcVoltage_2[30] ), 
        .\abcVoltage_2[31] (\abcVoltage_2[31] ), .\Min_out1[31] (Min_out1[31]), 
        .\Min_out1[19] (Min_out1[19]), .\Min_out1[20] (Min_out1[20]), .\Min_out1[21] (Min_out1[21]), 
        .\Gain1_mul_temp[9] (\Gain1_mul_temp[9] ), .\Min_out1[9] (Min_out1[9]), 
        .\Min_out1[22] (Min_out1[22]), .\Min_out1[23] (Min_out1[23]), .\Min_out1[24] (Min_out1[24]), 
        .\Min_out1[25] (Min_out1[25]), .\Min_out1[26] (Min_out1[26]), .\Min_out1[27] (Min_out1[27]), 
        .\Min_out1[28] (Min_out1[28]), .\Gain1_mul_temp[10] (\Gain1_mul_temp[10] ), 
        .\Min_out1[10] (Min_out1[10]), .\Gain1_mul_temp[13] (\Gain1_mul_temp[13] ), 
        .\Min_out1[13] (Min_out1[13]), .\Gain1_mul_temp[7] (\Gain1_mul_temp[7] ), 
        .\Min_out1[7] (Min_out1[7]), .\Gain1_mul_temp[6] (\Gain1_mul_temp[6] ), 
        .\Min_out1[6] (Min_out1[6]), .\Gain1_mul_temp[8] (\Gain1_mul_temp[8] ), 
        .\Min_out1[8] (Min_out1[8]), .\abcVoltage_1[14] (\abcVoltage_1[14] ), 
        .\Min_out1[14] (Min_out1[14]), .\Min_out1[29] (Min_out1[29]), .\Min_out1[30] (Min_out1[30]), 
        .\Gain1_mul_temp[4] (\Gain1_mul_temp[4] ), .\Min_out1[4] (Min_out1[4]), 
        .\Min_out1[12] (Min_out1[12]), .\Gain1_mul_temp[11] (\Gain1_mul_temp[11] ), 
        .\Min_out1[11] (Min_out1[11])) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/Space_Vector_Modulation.v(67[7] 71[15])
    Max u_Max (.\abcVoltage_1[31] (\abcVoltage_1[31] ), .alphaVoltage({alphaVoltage}), 
        .GND_net(GND_net), .\Gain1_mul_temp[11] (\Gain1_mul_temp[11] ), 
        .\abcVoltage_2[11] (\abcVoltage_2[11] ), .\Max_out1[11] (Max_out1[11]), 
        .\abcVoltage_1[17] (\abcVoltage_1[17] ), .\abcVoltage_1[16] (\abcVoltage_1[16] ), 
        .\abcVoltage_1[30] (\abcVoltage_1[30] ), .\Gain1_mul_temp[12] (\Gain1_mul_temp[12] ), 
        .\abcVoltage_2[12] (\abcVoltage_2[12] ), .\Max_out1[12] (Max_out1[12]), 
        .\Gain1_mul_temp[10] (\Gain1_mul_temp[10] ), .\abcVoltage_2[10] (\abcVoltage_2[10] ), 
        .\Max_out1[10] (Max_out1[10]), .\Gain1_mul_temp[5] (\Gain1_mul_temp[5] ), 
        .\abcVoltage_2[5] (\abcVoltage_2[5] ), .\Max_out1[5] (Max_out1[5]), 
        .\Gain1_mul_temp[9] (\Gain1_mul_temp[9] ), .\abcVoltage_2[9] (\abcVoltage_2[9] ), 
        .\Max_out1[9] (Max_out1[9]), .\Gain1_mul_temp[13] (\Gain1_mul_temp[13] ), 
        .\abcVoltage_2[13] (\abcVoltage_2[13] ), .\Max_out1[13] (Max_out1[13]), 
        .\Gain1_mul_temp[8] (\Gain1_mul_temp[8] ), .\abcVoltage_2[8] (\abcVoltage_2[8] ), 
        .\Max_out1[8] (Max_out1[8]), .\Gain1_mul_temp[6] (\Gain1_mul_temp[6] ), 
        .\abcVoltage_2[6] (\abcVoltage_2[6] ), .\Max_out1[6] (Max_out1[6]), 
        .\Gain1_mul_temp[7] (\Gain1_mul_temp[7] ), .\abcVoltage_2[7] (\abcVoltage_2[7] ), 
        .\Max_out1[7] (Max_out1[7]), .\abcVoltage_2[1] (\abcVoltage_2[1] ), 
        .\Max_out1[1] (Max_out1[1]), .\abcVoltage_1[14] (\abcVoltage_1[14] ), 
        .\abcVoltage_2[14] (\abcVoltage_2[14] ), .\Max_out1[14] (Max_out1[14]), 
        .\abcVoltage_2[2] (\abcVoltage_2[2] ), .\Max_out1[2] (Max_out1[2]), 
        .\Gain1_mul_temp[4] (\Gain1_mul_temp[4] ), .\abcVoltage_2[4] (\abcVoltage_2[4] ), 
        .\Max_out1[4] (Max_out1[4]), .\Gain1_mul_temp[3] (\Gain1_mul_temp[3] ), 
        .\abcVoltage_2[3] (\abcVoltage_2[3] ), .\Max_out1[3] (Max_out1[3]), 
        .\abcVoltage_2[15] (\abcVoltage_2[15] ), .\Max_out1[15] (Max_out1[15]), 
        .\abcVoltage_2[16] (\abcVoltage_2[16] ), .\Max_out1[16] (Max_out1[16]), 
        .\abcVoltage_2[17] (\abcVoltage_2[17] ), .\Max_out1[17] (Max_out1[17]), 
        .\abcVoltage_2[18] (\abcVoltage_2[18] ), .\Max_out1[18] (Max_out1[18]), 
        .\abcVoltage_2[31] (\abcVoltage_2[31] ), .\Max_out1[31] (Max_out1[31]), 
        .\abcVoltage_2[19] (\abcVoltage_2[19] ), .\Max_out1[19] (Max_out1[19]), 
        .\abcVoltage_2[20] (\abcVoltage_2[20] ), .\Max_out1[20] (Max_out1[20]), 
        .\abcVoltage_2[21] (\abcVoltage_2[21] ), .\Max_out1[21] (Max_out1[21]), 
        .\abcVoltage_2[22] (\abcVoltage_2[22] ), .\Max_out1[22] (Max_out1[22]), 
        .\abcVoltage_2[23] (\abcVoltage_2[23] ), .\Max_out1[23] (Max_out1[23]), 
        .\abcVoltage_2[24] (\abcVoltage_2[24] ), .\Max_out1[24] (Max_out1[24]), 
        .\abcVoltage_2[25] (\abcVoltage_2[25] ), .\Max_out1[25] (Max_out1[25]), 
        .\abcVoltage_2[26] (\abcVoltage_2[26] ), .\Max_out1[26] (Max_out1[26]), 
        .\abcVoltage_2[27] (\abcVoltage_2[27] ), .\Max_out1[27] (Max_out1[27]), 
        .\abcVoltage_2[28] (\abcVoltage_2[28] ), .\Max_out1[28] (Max_out1[28]), 
        .\abcVoltage_2[29] (\abcVoltage_2[29] ), .\Max_out1[29] (Max_out1[29]), 
        .\abcVoltage_2[30] (\abcVoltage_2[30] ), .\Max_out1[30] (Max_out1[30]), 
        .\abcVoltage_1[29] (\abcVoltage_1[29] ), .\abcVoltage_1[28] (\abcVoltage_1[28] ), 
        .\abcVoltage_1[27] (\abcVoltage_1[27] ), .\abcVoltage_1[26] (\abcVoltage_1[26] ), 
        .\abcVoltage_1[23] (\abcVoltage_1[23] ), .\abcVoltage_1[22] (\abcVoltage_1[22] ), 
        .\abcVoltage_1[18] (\abcVoltage_1[18] ), .\abcVoltage_1[15] (\abcVoltage_1[15] ), 
        .\Gain1_mul_temp[1] (\Gain1_mul_temp[1] ), .\Gain1_mul_temp[2] (\Gain1_mul_temp[2] ), 
        .\abcVoltage_1[21] (\abcVoltage_1[21] ), .\abcVoltage_1[20] (\abcVoltage_1[20] ), 
        .\abcVoltage_1[19] (\abcVoltage_1[19] ), .\abcVoltage_1[25] (\abcVoltage_1[25] ), 
        .\abcVoltage_1[24] (\abcVoltage_1[24] )) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/Space_Vector_Modulation.v(57[7] 61[15])
    VCC i1 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module Min
//

module Min (\abcVoltage_1[30] , alphaVoltage, GND_net, \Gain1_mul_temp[2] , 
            \Gain1_mul_temp[1] , \abcVoltage_1[26] , \abcVoltage_2[26] , 
            \abcVoltage_1[29] , \abcVoltage_2[29] , \abcVoltage_1[28] , 
            \abcVoltage_2[28] , \abcVoltage_1[27] , \abcVoltage_2[27] , 
            \abcVoltage_1[19] , \abcVoltage_2[19] , \abcVoltage_1[21] , 
            \abcVoltage_1[20] , \abcVoltage_2[20] , \abcVoltage_2[21] , 
            \abcVoltage_1[16] , \abcVoltage_1[15] , \abcVoltage_2[15] , 
            \abcVoltage_2[16] , \Gain1_mul_temp[3] , \abcVoltage_1[18] , 
            \abcVoltage_2[18] , \abcVoltage_1[17] , \abcVoltage_2[17] , 
            \abcVoltage_1[25] , \abcVoltage_1[23] , \abcVoltage_1[24] , 
            \abcVoltage_2[23] , \abcVoltage_2[24] , \abcVoltage_2[25] , 
            \abcVoltage_1[22] , \Gain1_mul_temp[12] , \abcVoltage_2[12] , 
            \abcVoltage_2[22] , \abcVoltage_1[31] , \abcVoltage_2[11] , 
            \abcVoltage_2[8] , \abcVoltage_2[6] , \abcVoltage_2[7] , \abcVoltage_2[3] , 
            \abcVoltage_2[1] , \Min_out1[1] , \abcVoltage_2[2] , \Min_out1[2] , 
            \Min_out1[3] , \abcVoltage_2[10] , \abcVoltage_2[5] , \abcVoltage_2[9] , 
            \abcVoltage_2[4] , \abcVoltage_2[13] , \Gain1_mul_temp[5] , 
            \abcVoltage_2[14] , \Min_out1[5] , \Min_out1[15] , \Min_out1[16] , 
            \Min_out1[17] , \Min_out1[18] , \abcVoltage_2[30] , \abcVoltage_2[31] , 
            \Min_out1[31] , \Min_out1[19] , \Min_out1[20] , \Min_out1[21] , 
            \Gain1_mul_temp[9] , \Min_out1[9] , \Min_out1[22] , \Min_out1[23] , 
            \Min_out1[24] , \Min_out1[25] , \Min_out1[26] , \Min_out1[27] , 
            \Min_out1[28] , \Gain1_mul_temp[10] , \Min_out1[10] , \Gain1_mul_temp[13] , 
            \Min_out1[13] , \Gain1_mul_temp[7] , \Min_out1[7] , \Gain1_mul_temp[6] , 
            \Min_out1[6] , \Gain1_mul_temp[8] , \Min_out1[8] , \abcVoltage_1[14] , 
            \Min_out1[14] , \Min_out1[29] , \Min_out1[30] , \Gain1_mul_temp[4] , 
            \Min_out1[4] , \Min_out1[12] , \Gain1_mul_temp[11] , \Min_out1[11] ) /* synthesis syn_module_defined=1 */ ;
    input \abcVoltage_1[30] ;
    input [15:0]alphaVoltage;
    input GND_net;
    input \Gain1_mul_temp[2] ;
    input \Gain1_mul_temp[1] ;
    input \abcVoltage_1[26] ;
    input \abcVoltage_2[26] ;
    input \abcVoltage_1[29] ;
    input \abcVoltage_2[29] ;
    input \abcVoltage_1[28] ;
    input \abcVoltage_2[28] ;
    input \abcVoltage_1[27] ;
    input \abcVoltage_2[27] ;
    input \abcVoltage_1[19] ;
    input \abcVoltage_2[19] ;
    input \abcVoltage_1[21] ;
    input \abcVoltage_1[20] ;
    input \abcVoltage_2[20] ;
    input \abcVoltage_2[21] ;
    input \abcVoltage_1[16] ;
    input \abcVoltage_1[15] ;
    input \abcVoltage_2[15] ;
    input \abcVoltage_2[16] ;
    input \Gain1_mul_temp[3] ;
    input \abcVoltage_1[18] ;
    input \abcVoltage_2[18] ;
    input \abcVoltage_1[17] ;
    input \abcVoltage_2[17] ;
    input \abcVoltage_1[25] ;
    input \abcVoltage_1[23] ;
    input \abcVoltage_1[24] ;
    input \abcVoltage_2[23] ;
    input \abcVoltage_2[24] ;
    input \abcVoltage_2[25] ;
    input \abcVoltage_1[22] ;
    input \Gain1_mul_temp[12] ;
    input \abcVoltage_2[12] ;
    input \abcVoltage_2[22] ;
    input \abcVoltage_1[31] ;
    input \abcVoltage_2[11] ;
    input \abcVoltage_2[8] ;
    input \abcVoltage_2[6] ;
    input \abcVoltage_2[7] ;
    input \abcVoltage_2[3] ;
    input \abcVoltage_2[1] ;
    output \Min_out1[1] ;
    input \abcVoltage_2[2] ;
    output \Min_out1[2] ;
    output \Min_out1[3] ;
    input \abcVoltage_2[10] ;
    input \abcVoltage_2[5] ;
    input \abcVoltage_2[9] ;
    input \abcVoltage_2[4] ;
    input \abcVoltage_2[13] ;
    input \Gain1_mul_temp[5] ;
    input \abcVoltage_2[14] ;
    output \Min_out1[5] ;
    output \Min_out1[15] ;
    output \Min_out1[16] ;
    output \Min_out1[17] ;
    output \Min_out1[18] ;
    input \abcVoltage_2[30] ;
    input \abcVoltage_2[31] ;
    output \Min_out1[31] ;
    output \Min_out1[19] ;
    output \Min_out1[20] ;
    output \Min_out1[21] ;
    input \Gain1_mul_temp[9] ;
    output \Min_out1[9] ;
    output \Min_out1[22] ;
    output \Min_out1[23] ;
    output \Min_out1[24] ;
    output \Min_out1[25] ;
    output \Min_out1[26] ;
    output \Min_out1[27] ;
    output \Min_out1[28] ;
    input \Gain1_mul_temp[10] ;
    output \Min_out1[10] ;
    input \Gain1_mul_temp[13] ;
    output \Min_out1[13] ;
    input \Gain1_mul_temp[7] ;
    output \Min_out1[7] ;
    input \Gain1_mul_temp[6] ;
    output \Min_out1[6] ;
    input \Gain1_mul_temp[8] ;
    output \Min_out1[8] ;
    input \abcVoltage_1[14] ;
    output \Min_out1[14] ;
    output \Min_out1[29] ;
    output \Min_out1[30] ;
    input \Gain1_mul_temp[4] ;
    output \Min_out1[4] ;
    output \Min_out1[12] ;
    input \Gain1_mul_temp[11] ;
    output \Min_out1[11] ;
    
    
    wire Min_stage1_val_0__31__N_337;
    wire [31:0]\Min_stage1_val[0] ;   // ../../hdlcoderFocCurrentFixptHdl/Min.v(35[22:36])
    
    wire n53, n59, n57, n55, n39, n41, n43, n31, n33, n37, 
        n35, n47, n49, n51, n25, n45, n59_adj_2192, n53_adj_2193, 
        n55_adj_2194, n47_adj_2195, n49_adj_2196, n51_adj_2197, n37_adj_2198, 
        n39_adj_2199, n41_adj_2200, n43_adj_2201, n45_adj_2202, n57_adj_2203, 
        n21649, n21736, n21836, n21832, n21651, n34, n21952, n21953, 
        n40, n21904, n42, n21691, n38, n36, n46, n21499, n22043, 
        n22044, n22018, n21906, n21919, n21986, n21921, n23, n21616, 
        n20, n21, n19, n11, n21618, n27, n21573, n21932, n29, 
        n17, n15, n13, n21606, n14, n12, n32, n9, n21634, 
        n21810, n21806, n22015, out0_31__N_336, n21892, n22033, 
        n21575, n21934, n18, n10, n26, n21567, n21995, n21996, 
        n8, n21870, n21871, n21742, n21922, n21705, n21947, n21744, 
        n21944, n21703, n6, n21950, n21951, n21600, n21592, n21993, 
        n21693, n22049, n22050, n22032, n22051, n22029, n21699, 
        n22059, n21710;
    
    SB_LUT4 in0_1_31__I_0_9_i31_3_lut (.I0(\abcVoltage_1[30] ), .I1(alphaVoltage[15]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [30]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13126_2_lut (.I0(\Gain1_mul_temp[2] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(GND_net), .I3(GND_net), .O(\Min_stage1_val[0] [2]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam i13126_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13125_2_lut (.I0(\Gain1_mul_temp[1] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(GND_net), .I3(GND_net), .O(\Min_stage1_val[0] [1]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam i13125_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 in0_1_31__I_0_9_i27_3_lut (.I0(\abcVoltage_1[26] ), .I1(alphaVoltage[11]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [26]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i53_2_lut (.I0(\Min_stage1_val[0] [26]), .I1(\abcVoltage_2[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i53_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i30_3_lut (.I0(\abcVoltage_1[29] ), .I1(alphaVoltage[14]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [29]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i59_2_lut (.I0(\Min_stage1_val[0] [29]), .I1(\abcVoltage_2[29] ), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i59_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i29_3_lut (.I0(\abcVoltage_1[28] ), .I1(alphaVoltage[13]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [28]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i57_2_lut (.I0(\Min_stage1_val[0] [28]), .I1(\abcVoltage_2[28] ), 
            .I2(GND_net), .I3(GND_net), .O(n57));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i57_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i28_3_lut (.I0(\abcVoltage_1[27] ), .I1(alphaVoltage[12]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [27]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i55_2_lut (.I0(\Min_stage1_val[0] [27]), .I1(\abcVoltage_2[27] ), 
            .I2(GND_net), .I3(GND_net), .O(n55));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i55_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i20_3_lut (.I0(\abcVoltage_1[19] ), .I1(alphaVoltage[4]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [19]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i39_2_lut (.I0(\Min_stage1_val[0] [19]), .I1(\abcVoltage_2[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i22_3_lut (.I0(\abcVoltage_1[21] ), .I1(alphaVoltage[6]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [21]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_9_i21_3_lut (.I0(\abcVoltage_1[20] ), .I1(alphaVoltage[5]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [20]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i41_2_lut (.I0(\Min_stage1_val[0] [20]), .I1(\abcVoltage_2[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_2_31__I_0_i43_2_lut (.I0(\Min_stage1_val[0] [21]), .I1(\abcVoltage_2[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i17_3_lut (.I0(\abcVoltage_1[16] ), .I1(alphaVoltage[1]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [16]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_9_i16_3_lut (.I0(\abcVoltage_1[15] ), .I1(alphaVoltage[0]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [15]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i31_2_lut (.I0(\Min_stage1_val[0] [15]), .I1(\abcVoltage_2[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_2_31__I_0_i33_2_lut (.I0(\Min_stage1_val[0] [16]), .I1(\abcVoltage_2[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13127_2_lut (.I0(\Gain1_mul_temp[3] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(GND_net), .I3(GND_net), .O(\Min_stage1_val[0] [3]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam i13127_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 in0_1_31__I_0_9_i19_3_lut (.I0(\abcVoltage_1[18] ), .I1(alphaVoltage[3]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [18]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i37_2_lut (.I0(\Min_stage1_val[0] [18]), .I1(\abcVoltage_2[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i18_3_lut (.I0(\abcVoltage_1[17] ), .I1(alphaVoltage[2]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [17]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i35_2_lut (.I0(\Min_stage1_val[0] [17]), .I1(\abcVoltage_2[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i26_3_lut (.I0(\abcVoltage_1[25] ), .I1(alphaVoltage[10]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [25]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_9_i24_3_lut (.I0(\abcVoltage_1[23] ), .I1(alphaVoltage[8]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [23]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_9_i25_3_lut (.I0(\abcVoltage_1[24] ), .I1(alphaVoltage[9]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [24]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i47_2_lut (.I0(\Min_stage1_val[0] [23]), .I1(\abcVoltage_2[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i47_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_2_31__I_0_i49_2_lut (.I0(\Min_stage1_val[0] [24]), .I1(\abcVoltage_2[24] ), 
            .I2(GND_net), .I3(GND_net), .O(n49));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i49_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_2_31__I_0_i51_2_lut (.I0(\Min_stage1_val[0] [25]), .I1(\abcVoltage_2[25] ), 
            .I2(GND_net), .I3(GND_net), .O(n51));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i51_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_9_i23_3_lut (.I0(\abcVoltage_1[22] ), .I1(alphaVoltage[7]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [22]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i25_2_lut_3_lut (.I0(\Gain1_mul_temp[12] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[12] ), .I3(GND_net), .O(n25));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i25_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i45_2_lut (.I0(\Min_stage1_val[0] [22]), .I1(\abcVoltage_2[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i59_2_lut (.I0(alphaVoltage[14]), .I1(\abcVoltage_1[29] ), 
            .I2(GND_net), .I3(GND_net), .O(n59_adj_2192));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i59_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i53_2_lut (.I0(alphaVoltage[11]), .I1(\abcVoltage_1[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_2193));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i53_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i55_2_lut (.I0(alphaVoltage[12]), .I1(\abcVoltage_1[27] ), 
            .I2(GND_net), .I3(GND_net), .O(n55_adj_2194));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i55_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i47_2_lut (.I0(alphaVoltage[8]), .I1(\abcVoltage_1[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_2195));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i47_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i49_2_lut (.I0(alphaVoltage[9]), .I1(\abcVoltage_1[24] ), 
            .I2(GND_net), .I3(GND_net), .O(n49_adj_2196));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i49_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i51_2_lut (.I0(alphaVoltage[10]), .I1(\abcVoltage_1[25] ), 
            .I2(GND_net), .I3(GND_net), .O(n51_adj_2197));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i51_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i37_2_lut (.I0(alphaVoltage[3]), .I1(\abcVoltage_1[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_2198));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i39_2_lut (.I0(alphaVoltage[4]), .I1(\abcVoltage_1[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_2199));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i41_2_lut (.I0(alphaVoltage[5]), .I1(\abcVoltage_1[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_2200));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i43_2_lut (.I0(alphaVoltage[6]), .I1(\abcVoltage_1[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_2201));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i45_2_lut (.I0(alphaVoltage[7]), .I1(\abcVoltage_1[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_2202));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i57_2_lut (.I0(alphaVoltage[13]), .I1(\abcVoltage_1[28] ), 
            .I2(GND_net), .I3(GND_net), .O(n57_adj_2203));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i57_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16637_4_lut (.I0(n57_adj_2203), .I1(n45_adj_2202), .I2(n43_adj_2201), 
            .I3(n41_adj_2200), .O(n21649));
    defparam i16637_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16724_4_lut (.I0(n39_adj_2199), .I1(n37_adj_2198), .I2(alphaVoltage[2]), 
            .I3(\abcVoltage_1[17] ), .O(n21736));
    defparam i16724_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i16824_4_lut (.I0(n45_adj_2202), .I1(n43_adj_2201), .I2(n41_adj_2200), 
            .I3(n21736), .O(n21836));
    defparam i16824_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i16820_4_lut (.I0(n51_adj_2197), .I1(n49_adj_2196), .I2(n47_adj_2195), 
            .I3(n21836), .O(n21832));
    defparam i16820_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i16639_4_lut (.I0(n57_adj_2203), .I1(n55_adj_2194), .I2(n53_adj_2193), 
            .I3(n21832), .O(n21651));
    defparam i16639_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 in0_1_31__I_0_i34_4_lut (.I0(\abcVoltage_1[15] ), .I1(\abcVoltage_1[16] ), 
            .I2(alphaVoltage[1]), .I3(alphaVoltage[0]), .O(n34));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i34_4_lut.LUT_INIT = 16'h8ecf;
    SB_LUT4 i16940_3_lut (.I0(n34), .I1(\abcVoltage_1[28] ), .I2(n57_adj_2203), 
            .I3(GND_net), .O(n21952));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i16940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16941_3_lut (.I0(n21952), .I1(\abcVoltage_1[29] ), .I2(n59_adj_2192), 
            .I3(GND_net), .O(n21953));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i16941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i40_3_lut (.I0(\abcVoltage_1[20] ), .I1(\abcVoltage_1[21] ), 
            .I2(n43_adj_2201), .I3(GND_net), .O(n40));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16892_4_lut (.I0(alphaVoltage[15]), .I1(n59_adj_2192), .I2(\abcVoltage_1[30] ), 
            .I3(n21649), .O(n21904));
    defparam i16892_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 in0_1_31__I_0_i42_3_lut (.I0(n40), .I1(\abcVoltage_1[22] ), 
            .I2(n45_adj_2202), .I3(GND_net), .O(n42));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16679_3_lut (.I0(n21953), .I1(\abcVoltage_1[30] ), .I2(alphaVoltage[15]), 
            .I3(GND_net), .O(n21691));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i16679_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 in0_1_31__I_0_i38_3_lut (.I0(\abcVoltage_1[19] ), .I1(\abcVoltage_1[23] ), 
            .I2(n47_adj_2195), .I3(GND_net), .O(n38));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i36_3_lut (.I0(\abcVoltage_1[17] ), .I1(\abcVoltage_1[18] ), 
            .I2(n37_adj_2198), .I3(GND_net), .O(n36));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i46_3_lut (.I0(n38), .I1(\abcVoltage_1[24] ), 
            .I2(n49_adj_2196), .I3(GND_net), .O(n46));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i46_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17031_4_lut (.I0(n46), .I1(n36), .I2(n49_adj_2196), .I3(n21499), 
            .O(n22043));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i17031_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i17032_3_lut (.I0(n22043), .I1(\abcVoltage_1[25] ), .I2(n51_adj_2197), 
            .I3(GND_net), .O(n22044));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i17032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17006_3_lut (.I0(n22044), .I1(\abcVoltage_1[26] ), .I2(n53_adj_2193), 
            .I3(GND_net), .O(n22018));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i17006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16894_4_lut (.I0(alphaVoltage[15]), .I1(n59_adj_2192), .I2(\abcVoltage_1[30] ), 
            .I3(n21651), .O(n21906));
    defparam i16894_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i16907_3_lut (.I0(n21691), .I1(n42), .I2(n21904), .I3(GND_net), 
            .O(n21919));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i16907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16974_3_lut (.I0(n22018), .I1(\abcVoltage_1[27] ), .I2(n55_adj_2194), 
            .I3(GND_net), .O(n21986));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i16974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16909_3_lut (.I0(n21986), .I1(n21919), .I2(n21906), .I3(GND_net), 
            .O(n21921));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam i16909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i64_3_lut (.I0(n21921), .I1(alphaVoltage[15]), 
            .I2(\abcVoltage_1[31] ), .I3(GND_net), .O(Min_stage1_val_0__31__N_337));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[31:47])
    defparam in0_1_31__I_0_i64_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16604_2_lut (.I0(n25), .I1(n23), .I2(GND_net), .I3(GND_net), 
            .O(n21616));
    defparam i16604_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 in0_2_31__I_0_i20_3_lut (.I0(\abcVoltage_2[11] ), .I1(\abcVoltage_2[12] ), 
            .I2(n25), .I3(GND_net), .O(n20));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16606_4_lut (.I0(n23), .I1(n21), .I2(n19), .I3(n11), .O(n21618));
    defparam i16606_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16561_4_lut (.I0(n45), .I1(n27), .I2(n25), .I3(n21618), 
            .O(n21573));
    defparam i16561_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16920_4_lut (.I0(n51), .I1(n49), .I2(n47), .I3(n21573), 
            .O(n21932));
    defparam i16920_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16594_4_lut (.I0(n29), .I1(n17), .I2(n15), .I3(n13), .O(n21606));
    defparam i16594_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 in0_2_31__I_0_i14_3_lut (.I0(\abcVoltage_2[8] ), .I1(\abcVoltage_2[17] ), 
            .I2(n35), .I3(GND_net), .O(n14));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i12_3_lut (.I0(\abcVoltage_2[6] ), .I1(\abcVoltage_2[7] ), 
            .I2(n15), .I3(GND_net), .O(n12));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i32_3_lut (.I0(n14), .I1(\abcVoltage_2[18] ), 
            .I2(n37), .I3(GND_net), .O(n32));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16622_3_lut (.I0(n9), .I1(\Min_stage1_val[0] [3]), .I2(\abcVoltage_2[3] ), 
            .I3(GND_net), .O(n21634));
    defparam i16622_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i16798_4_lut (.I0(n15), .I1(n13), .I2(n11), .I3(n21634), 
            .O(n21810));
    defparam i16798_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i16794_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n21810), 
            .O(n21806));
    defparam i16794_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i17003_4_lut (.I0(n27), .I1(n25), .I2(n23), .I3(n21806), 
            .O(n22015));
    defparam i17003_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 in0_2_31__I_0_8_i2_3_lut (.I0(\abcVoltage_2[1] ), .I1(\Min_stage1_val[0] [1]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[1] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i3_3_lut (.I0(\abcVoltage_2[2] ), .I1(\Min_stage1_val[0] [2]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[2] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i4_3_lut (.I0(\abcVoltage_2[3] ), .I1(\Min_stage1_val[0] [3]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[3] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16880_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n22015), 
            .O(n21892));
    defparam i16880_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i17021_4_lut (.I0(n39), .I1(n37), .I2(n35), .I3(n21892), 
            .O(n22033));
    defparam i17021_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16563_4_lut (.I0(n45), .I1(n43), .I2(n41), .I3(n22033), 
            .O(n21575));
    defparam i16563_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16922_4_lut (.I0(n51), .I1(n49), .I2(n47), .I3(n21575), 
            .O(n21934));
    defparam i16922_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 in0_2_31__I_0_i18_3_lut (.I0(\abcVoltage_2[10] ), .I1(\abcVoltage_2[22] ), 
            .I2(n45), .I3(GND_net), .O(n18));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i10_3_lut (.I0(\abcVoltage_2[5] ), .I1(\abcVoltage_2[9] ), 
            .I2(n19), .I3(GND_net), .O(n10));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i26_3_lut (.I0(n18), .I1(\abcVoltage_2[23] ), 
            .I2(n47), .I3(GND_net), .O(n26));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16983_4_lut (.I0(n26), .I1(n10), .I2(n47), .I3(n21567), 
            .O(n21995));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16983_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i16984_3_lut (.I0(n21995), .I1(\abcVoltage_2[24] ), .I2(n49), 
            .I3(GND_net), .O(n21996));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i8_3_lut (.I0(\abcVoltage_2[3] ), .I1(\abcVoltage_2[4] ), 
            .I2(n9), .I3(GND_net), .O(n8));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16858_3_lut (.I0(n8), .I1(\abcVoltage_2[27] ), .I2(n55), 
            .I3(GND_net), .O(n21870));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16859_3_lut (.I0(n21870), .I1(\abcVoltage_2[28] ), .I2(n57), 
            .I3(GND_net), .O(n21871));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16730_4_lut (.I0(n57), .I1(n55), .I2(n27), .I3(n21616), 
            .O(n21742));
    defparam i16730_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i16910_3_lut (.I0(n20), .I1(\abcVoltage_2[13] ), .I2(n27), 
            .I3(GND_net), .O(n21922));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16693_3_lut (.I0(n21871), .I1(\abcVoltage_2[29] ), .I2(n59), 
            .I3(GND_net), .O(n21705));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16935_3_lut (.I0(n21996), .I1(\abcVoltage_2[25] ), .I2(n51), 
            .I3(GND_net), .O(n21947));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16732_4_lut (.I0(n57), .I1(n55), .I2(n53), .I3(n21932), 
            .O(n21744));
    defparam i16732_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 in0_2_31__I_0_i11_2_lut_3_lut (.I0(\Gain1_mul_temp[5] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[5] ), .I3(GND_net), .O(n11));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i11_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i16932_4_lut (.I0(n21705), .I1(n21922), .I2(n59), .I3(n21742), 
            .O(n21944));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16932_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i16691_3_lut (.I0(n21947), .I1(\abcVoltage_2[26] ), .I2(n53), 
            .I3(GND_net), .O(n21703));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i6_4_lut (.I0(\Min_stage1_val[0] [1]), .I1(\abcVoltage_2[2] ), 
            .I2(\Min_stage1_val[0] [2]), .I3(\abcVoltage_2[1] ), .O(n6));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam in0_2_31__I_0_i6_4_lut.LUT_INIT = 16'hcf4d;
    SB_LUT4 i16938_3_lut (.I0(n6), .I1(\abcVoltage_2[14] ), .I2(n29), 
            .I3(GND_net), .O(n21950));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i6_3_lut_4_lut (.I0(\Gain1_mul_temp[5] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[5] ), .O(\Min_out1[5] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i6_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i16939_3_lut (.I0(n21950), .I1(\abcVoltage_2[15] ), .I2(n31), 
            .I3(GND_net), .O(n21951));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16588_4_lut (.I0(n35), .I1(n33), .I2(n31), .I3(n21606), 
            .O(n21600));
    defparam i16588_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16981_4_lut (.I0(n32), .I1(n12), .I2(n37), .I3(n21592), 
            .O(n21993));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16981_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i16681_3_lut (.I0(n21951), .I1(\abcVoltage_2[16] ), .I2(n33), 
            .I3(GND_net), .O(n21693));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i16_3_lut (.I0(\abcVoltage_2[15] ), .I1(\Min_stage1_val[0] [15]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[15] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i17_3_lut (.I0(\abcVoltage_2[16] ), .I1(\Min_stage1_val[0] [16]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[16] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17037_4_lut (.I0(n21693), .I1(n21993), .I2(n37), .I3(n21600), 
            .O(n22049));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i17037_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i17038_3_lut (.I0(n22049), .I1(\abcVoltage_2[19] ), .I2(n39), 
            .I3(GND_net), .O(n22050));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i17038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17020_3_lut (.I0(n22050), .I1(\abcVoltage_2[20] ), .I2(n41), 
            .I3(GND_net), .O(n22032));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i17020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17039_4_lut (.I0(n57), .I1(n55), .I2(n53), .I3(n21934), 
            .O(n22051));
    defparam i17039_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17017_4_lut (.I0(n21703), .I1(n21944), .I2(n59), .I3(n21744), 
            .O(n22029));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i17017_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 in0_2_31__I_0_8_i18_3_lut (.I0(\abcVoltage_2[17] ), .I1(\Min_stage1_val[0] [17]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[17] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i19_3_lut (.I0(\abcVoltage_2[18] ), .I1(\Min_stage1_val[0] [18]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[18] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16687_3_lut (.I0(n22032), .I1(\abcVoltage_2[21] ), .I2(n43), 
            .I3(GND_net), .O(n21699));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17047_4_lut (.I0(n21699), .I1(n22029), .I2(n59), .I3(n22051), 
            .O(n22059));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i17047_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16698_3_lut (.I0(n22059), .I1(\abcVoltage_2[30] ), .I2(\Min_stage1_val[0] [30]), 
            .I3(GND_net), .O(n21710));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16698_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16699_3_lut (.I0(n21710), .I1(\Min_stage1_val[0] [31]), .I2(\abcVoltage_2[31] ), 
            .I3(GND_net), .O(out0_31__N_336));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[28:66])
    defparam i16699_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 in0_1_31__I_0_9_i32_3_lut (.I0(\abcVoltage_1[31] ), .I1(alphaVoltage[15]), 
            .I2(Min_stage1_val_0__31__N_337), .I3(GND_net), .O(\Min_stage1_val[0] [31]));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_1_31__I_0_9_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i32_3_lut (.I0(\abcVoltage_2[31] ), .I1(\Min_stage1_val[0] [31]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[31] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i20_3_lut (.I0(\abcVoltage_2[19] ), .I1(\Min_stage1_val[0] [19]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[19] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i21_3_lut (.I0(\abcVoltage_2[20] ), .I1(\Min_stage1_val[0] [20]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[20] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i22_3_lut (.I0(\abcVoltage_2[21] ), .I1(\Min_stage1_val[0] [21]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[21] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i19_2_lut_3_lut (.I0(\Gain1_mul_temp[9] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[9] ), .I3(GND_net), .O(n19));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i19_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i10_3_lut_4_lut (.I0(\Gain1_mul_temp[9] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[9] ), .O(\Min_out1[9] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i10_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_8_i23_3_lut (.I0(\abcVoltage_2[22] ), .I1(\Min_stage1_val[0] [22]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[22] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i24_3_lut (.I0(\abcVoltage_2[23] ), .I1(\Min_stage1_val[0] [23]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[23] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i25_3_lut (.I0(\abcVoltage_2[24] ), .I1(\Min_stage1_val[0] [24]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[24] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i26_3_lut (.I0(\abcVoltage_2[25] ), .I1(\Min_stage1_val[0] [25]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[25] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i27_3_lut (.I0(\abcVoltage_2[26] ), .I1(\Min_stage1_val[0] [26]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[26] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i28_3_lut (.I0(\abcVoltage_2[27] ), .I1(\Min_stage1_val[0] [27]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[27] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i29_3_lut (.I0(\abcVoltage_2[28] ), .I1(\Min_stage1_val[0] [28]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[28] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i21_2_lut_3_lut (.I0(\Gain1_mul_temp[10] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[10] ), .I3(GND_net), .O(n21));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i21_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i11_3_lut_4_lut (.I0(\Gain1_mul_temp[10] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[10] ), .O(\Min_out1[10] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i11_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_8_i14_3_lut_4_lut (.I0(\Gain1_mul_temp[13] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[13] ), .O(\Min_out1[13] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i14_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i27_2_lut_3_lut (.I0(\Gain1_mul_temp[13] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[13] ), .I3(GND_net), .O(n27));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i27_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i15_2_lut_3_lut (.I0(\Gain1_mul_temp[7] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[7] ), .I3(GND_net), .O(n15));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i15_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i8_3_lut_4_lut (.I0(\Gain1_mul_temp[7] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[7] ), .O(\Min_out1[7] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i8_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i13_2_lut_3_lut (.I0(\Gain1_mul_temp[6] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[6] ), .I3(GND_net), .O(n13));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i13_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i7_3_lut_4_lut (.I0(\Gain1_mul_temp[6] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[6] ), .O(\Min_out1[6] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i7_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i17_2_lut_3_lut (.I0(\Gain1_mul_temp[8] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[8] ), .I3(GND_net), .O(n17));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i17_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i9_3_lut_4_lut (.I0(\Gain1_mul_temp[8] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[8] ), .O(\Min_out1[8] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i9_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_8_i15_3_lut_4_lut (.I0(\abcVoltage_1[14] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[14] ), .O(\Min_out1[14] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i29_2_lut_3_lut (.I0(\abcVoltage_1[14] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[14] ), .I3(GND_net), .O(n29));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i29_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i30_3_lut (.I0(\abcVoltage_2[29] ), .I1(\Min_stage1_val[0] [29]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[29] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_8_i31_3_lut (.I0(\abcVoltage_2[30] ), .I1(\Min_stage1_val[0] [30]), 
            .I2(out0_31__N_336), .I3(GND_net), .O(\Min_out1[30] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(52[27] 53[33])
    defparam in0_2_31__I_0_8_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i9_2_lut_3_lut (.I0(\Gain1_mul_temp[4] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[4] ), .I3(GND_net), .O(n9));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i9_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i5_3_lut_4_lut (.I0(\Gain1_mul_temp[4] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[4] ), .O(\Min_out1[4] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i5_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_8_i13_3_lut_4_lut (.I0(\Gain1_mul_temp[12] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[12] ), .O(\Min_out1[12] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i13_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i23_2_lut_3_lut (.I0(\Gain1_mul_temp[11] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(\abcVoltage_2[11] ), .I3(GND_net), .O(n23));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_i23_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_8_i12_3_lut_4_lut (.I0(\Gain1_mul_temp[11] ), .I1(Min_stage1_val_0__31__N_337), 
            .I2(out0_31__N_336), .I3(\abcVoltage_2[11] ), .O(\Min_out1[11] ));   // ../../hdlcoderFocCurrentFixptHdl/Min.v(45[30] 46[22])
    defparam in0_2_31__I_0_8_i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i16555_2_lut_3_lut (.I0(\Min_stage1_val[0] [22]), .I1(\abcVoltage_2[22] ), 
            .I2(n21), .I3(GND_net), .O(n21567));
    defparam i16555_2_lut_3_lut.LUT_INIT = 16'hf6f6;
    SB_LUT4 i16580_2_lut_3_lut (.I0(\Min_stage1_val[0] [17]), .I1(\abcVoltage_2[17] ), 
            .I2(n17), .I3(GND_net), .O(n21592));
    defparam i16580_2_lut_3_lut.LUT_INIT = 16'hf6f6;
    SB_LUT4 i16493_2_lut_4_lut (.I0(alphaVoltage[8]), .I1(\abcVoltage_1[23] ), 
            .I2(alphaVoltage[4]), .I3(\abcVoltage_1[19] ), .O(n21499));
    defparam i16493_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    
endmodule
//
// Verilog Description of module Max
//

module Max (\abcVoltage_1[31] , alphaVoltage, GND_net, \Gain1_mul_temp[11] , 
            \abcVoltage_2[11] , \Max_out1[11] , \abcVoltage_1[17] , \abcVoltage_1[16] , 
            \abcVoltage_1[30] , \Gain1_mul_temp[12] , \abcVoltage_2[12] , 
            \Max_out1[12] , \Gain1_mul_temp[10] , \abcVoltage_2[10] , 
            \Max_out1[10] , \Gain1_mul_temp[5] , \abcVoltage_2[5] , \Max_out1[5] , 
            \Gain1_mul_temp[9] , \abcVoltage_2[9] , \Max_out1[9] , \Gain1_mul_temp[13] , 
            \abcVoltage_2[13] , \Max_out1[13] , \Gain1_mul_temp[8] , \abcVoltage_2[8] , 
            \Max_out1[8] , \Gain1_mul_temp[6] , \abcVoltage_2[6] , \Max_out1[6] , 
            \Gain1_mul_temp[7] , \abcVoltage_2[7] , \Max_out1[7] , \abcVoltage_2[1] , 
            \Max_out1[1] , \abcVoltage_1[14] , \abcVoltage_2[14] , \Max_out1[14] , 
            \abcVoltage_2[2] , \Max_out1[2] , \Gain1_mul_temp[4] , \abcVoltage_2[4] , 
            \Max_out1[4] , \Gain1_mul_temp[3] , \abcVoltage_2[3] , \Max_out1[3] , 
            \abcVoltage_2[15] , \Max_out1[15] , \abcVoltage_2[16] , \Max_out1[16] , 
            \abcVoltage_2[17] , \Max_out1[17] , \abcVoltage_2[18] , \Max_out1[18] , 
            \abcVoltage_2[31] , \Max_out1[31] , \abcVoltage_2[19] , \Max_out1[19] , 
            \abcVoltage_2[20] , \Max_out1[20] , \abcVoltage_2[21] , \Max_out1[21] , 
            \abcVoltage_2[22] , \Max_out1[22] , \abcVoltage_2[23] , \Max_out1[23] , 
            \abcVoltage_2[24] , \Max_out1[24] , \abcVoltage_2[25] , \Max_out1[25] , 
            \abcVoltage_2[26] , \Max_out1[26] , \abcVoltage_2[27] , \Max_out1[27] , 
            \abcVoltage_2[28] , \Max_out1[28] , \abcVoltage_2[29] , \Max_out1[29] , 
            \abcVoltage_2[30] , \Max_out1[30] , \abcVoltage_1[29] , \abcVoltage_1[28] , 
            \abcVoltage_1[27] , \abcVoltage_1[26] , \abcVoltage_1[23] , 
            \abcVoltage_1[22] , \abcVoltage_1[18] , \abcVoltage_1[15] , 
            \Gain1_mul_temp[1] , \Gain1_mul_temp[2] , \abcVoltage_1[21] , 
            \abcVoltage_1[20] , \abcVoltage_1[19] , \abcVoltage_1[25] , 
            \abcVoltage_1[24] ) /* synthesis syn_module_defined=1 */ ;
    input \abcVoltage_1[31] ;
    input [15:0]alphaVoltage;
    input GND_net;
    input \Gain1_mul_temp[11] ;
    input \abcVoltage_2[11] ;
    output \Max_out1[11] ;
    input \abcVoltage_1[17] ;
    input \abcVoltage_1[16] ;
    input \abcVoltage_1[30] ;
    input \Gain1_mul_temp[12] ;
    input \abcVoltage_2[12] ;
    output \Max_out1[12] ;
    input \Gain1_mul_temp[10] ;
    input \abcVoltage_2[10] ;
    output \Max_out1[10] ;
    input \Gain1_mul_temp[5] ;
    input \abcVoltage_2[5] ;
    output \Max_out1[5] ;
    input \Gain1_mul_temp[9] ;
    input \abcVoltage_2[9] ;
    output \Max_out1[9] ;
    input \Gain1_mul_temp[13] ;
    input \abcVoltage_2[13] ;
    output \Max_out1[13] ;
    input \Gain1_mul_temp[8] ;
    input \abcVoltage_2[8] ;
    output \Max_out1[8] ;
    input \Gain1_mul_temp[6] ;
    input \abcVoltage_2[6] ;
    output \Max_out1[6] ;
    input \Gain1_mul_temp[7] ;
    input \abcVoltage_2[7] ;
    output \Max_out1[7] ;
    input \abcVoltage_2[1] ;
    output \Max_out1[1] ;
    input \abcVoltage_1[14] ;
    input \abcVoltage_2[14] ;
    output \Max_out1[14] ;
    input \abcVoltage_2[2] ;
    output \Max_out1[2] ;
    input \Gain1_mul_temp[4] ;
    input \abcVoltage_2[4] ;
    output \Max_out1[4] ;
    input \Gain1_mul_temp[3] ;
    input \abcVoltage_2[3] ;
    output \Max_out1[3] ;
    input \abcVoltage_2[15] ;
    output \Max_out1[15] ;
    input \abcVoltage_2[16] ;
    output \Max_out1[16] ;
    input \abcVoltage_2[17] ;
    output \Max_out1[17] ;
    input \abcVoltage_2[18] ;
    output \Max_out1[18] ;
    input \abcVoltage_2[31] ;
    output \Max_out1[31] ;
    input \abcVoltage_2[19] ;
    output \Max_out1[19] ;
    input \abcVoltage_2[20] ;
    output \Max_out1[20] ;
    input \abcVoltage_2[21] ;
    output \Max_out1[21] ;
    input \abcVoltage_2[22] ;
    output \Max_out1[22] ;
    input \abcVoltage_2[23] ;
    output \Max_out1[23] ;
    input \abcVoltage_2[24] ;
    output \Max_out1[24] ;
    input \abcVoltage_2[25] ;
    output \Max_out1[25] ;
    input \abcVoltage_2[26] ;
    output \Max_out1[26] ;
    input \abcVoltage_2[27] ;
    output \Max_out1[27] ;
    input \abcVoltage_2[28] ;
    output \Max_out1[28] ;
    input \abcVoltage_2[29] ;
    output \Max_out1[29] ;
    input \abcVoltage_2[30] ;
    output \Max_out1[30] ;
    input \abcVoltage_1[29] ;
    input \abcVoltage_1[28] ;
    input \abcVoltage_1[27] ;
    input \abcVoltage_1[26] ;
    input \abcVoltage_1[23] ;
    input \abcVoltage_1[22] ;
    input \abcVoltage_1[18] ;
    input \abcVoltage_1[15] ;
    input \Gain1_mul_temp[1] ;
    input \Gain1_mul_temp[2] ;
    input \abcVoltage_1[21] ;
    input \abcVoltage_1[20] ;
    input \abcVoltage_1[19] ;
    input \abcVoltage_1[25] ;
    input \abcVoltage_1[24] ;
    
    
    wire Max_stage1_val_0__31__N_335;
    wire [31:0]\Max_stage1_val[0] ;   // ../../hdlcoderFocCurrentFixptHdl/Max.v(35[22:36])
    
    wire out0_31__N_334, n23, n21545, n34, n21914, n25, n21, n11, 
        n19, n27, n49, n22, n17, n13, n15, n29, n6, n16, 
        n9, n7, n47, n45, n33, n35, n37, n31, n38, n43, 
        n40, n56, n21842, n21912, n52, n21844, n39, n41, n43_adj_2183, 
        n51, n49_adj_2184, n51_adj_2185, n53, n45_adj_2186, n47_adj_2187, 
        n37_adj_2188, n41_adj_2189, n39_adj_2190, n21730, n21549, 
        n21926, n59, n57, n55, n36, n44, n21547, n22009, n22010, 
        n21961, n21660, n20038, n20044, n20050, n20056, n32, n21880, 
        n21881, n21647, n21515, n21768, n44_adj_2191, n21780, n21824, 
        n21882, n21638, n19887, n21497, n21632, n21938, n21820, 
        n22013, n21890, n21507, n21513, n21505, n21587, n21987, 
        n24, n42, n21956, n21957, n21868, n22041, n21681, n21509, 
        n21511, n21958, n21959, n21814, n22039, n21679, n22037, 
        n22072, n22060, n22087, n22088, n22086, n22074, n22075, 
        n22063;
    
    SB_LUT4 in0_1_31__I_0_i32_3_lut (.I0(\abcVoltage_1[31] ), .I1(alphaVoltage[15]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [31]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i12_3_lut_4_lut (.I0(\Gain1_mul_temp[11] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[11] ), .O(\Max_out1[11] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i23_2_lut_3_lut (.I0(\Gain1_mul_temp[11] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[11] ), .I3(GND_net), 
            .O(n23));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i23_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i16533_3_lut_4_lut (.I0(\abcVoltage_1[17] ), .I1(alphaVoltage[2]), 
            .I2(alphaVoltage[1]), .I3(\abcVoltage_1[16] ), .O(n21545));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16533_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 in0_0_31__I_0_i34_3_lut_3_lut (.I0(\abcVoltage_1[17] ), .I1(alphaVoltage[2]), 
            .I2(alphaVoltage[1]), .I3(GND_net), .O(n34));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i14905_3_lut_4_lut_4_lut (.I0(\abcVoltage_1[30] ), .I1(alphaVoltage[15]), 
            .I2(\abcVoltage_1[31] ), .I3(n21914), .O(Max_stage1_val_0__31__N_335));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i14905_3_lut_4_lut_4_lut.LUT_INIT = 16'hf170;
    SB_LUT4 Max_stage1_val_0__31__I_0_i25_2_lut_3_lut (.I0(\Gain1_mul_temp[12] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[12] ), .I3(GND_net), 
            .O(n25));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i25_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i13_3_lut_4_lut (.I0(\Gain1_mul_temp[12] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[12] ), .O(\Max_out1[12] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i13_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i11_3_lut_4_lut (.I0(\Gain1_mul_temp[10] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[10] ), .O(\Max_out1[10] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i11_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i21_2_lut_3_lut (.I0(\Gain1_mul_temp[10] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[10] ), .I3(GND_net), 
            .O(n21));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i21_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 Max_stage1_val_0__31__I_0_i11_2_lut_3_lut (.I0(\Gain1_mul_temp[5] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[5] ), .I3(GND_net), 
            .O(n11));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i11_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i6_3_lut_4_lut (.I0(\Gain1_mul_temp[5] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[5] ), .O(\Max_out1[5] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i6_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i10_3_lut_4_lut (.I0(\Gain1_mul_temp[9] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[9] ), .O(\Max_out1[9] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i10_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i19_2_lut_3_lut (.I0(\Gain1_mul_temp[9] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[9] ), .I3(GND_net), 
            .O(n19));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i19_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i14_3_lut_4_lut (.I0(\Gain1_mul_temp[13] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[13] ), .O(\Max_out1[13] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i14_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i27_2_lut_3_lut (.I0(\Gain1_mul_temp[13] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[13] ), .I3(GND_net), 
            .O(n27));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i27_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 Max_stage1_val_0__31__I_0_i22_3_lut_4_lut (.I0(\Gain1_mul_temp[13] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(n49), .I3(\Max_stage1_val[0] [24]), 
            .O(n22));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i22_3_lut_4_lut.LUT_INIT = 16'hf202;
    SB_LUT4 in0_2_31__I_0_i9_3_lut_4_lut (.I0(\Gain1_mul_temp[8] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[8] ), .O(\Max_out1[8] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i9_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i17_2_lut_3_lut (.I0(\Gain1_mul_temp[8] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[8] ), .I3(GND_net), 
            .O(n17));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i17_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 Max_stage1_val_0__31__I_0_i13_2_lut_3_lut (.I0(\Gain1_mul_temp[6] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[6] ), .I3(GND_net), 
            .O(n13));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i13_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i7_3_lut_4_lut (.I0(\Gain1_mul_temp[6] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[6] ), .O(\Max_out1[6] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i7_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i8_3_lut_4_lut (.I0(\Gain1_mul_temp[7] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[7] ), .O(\Max_out1[7] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i8_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i2_3_lut (.I0(\abcVoltage_2[1] ), .I1(\Max_stage1_val[0] [1]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[1] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i15_2_lut_3_lut (.I0(\Gain1_mul_temp[7] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[7] ), .I3(GND_net), 
            .O(n15));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i15_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 Max_stage1_val_0__31__I_0_i16_3_lut_4_lut (.I0(\abcVoltage_1[14] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(n29), .I3(n6), .O(n16));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i16_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i15_3_lut_4_lut (.I0(\abcVoltage_1[14] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[14] ), .O(\Max_out1[14] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i29_2_lut_3_lut (.I0(\abcVoltage_1[14] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[14] ), .I3(GND_net), 
            .O(n29));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i29_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i3_3_lut (.I0(\abcVoltage_2[2] ), .I1(\Max_stage1_val[0] [2]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[2] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i9_2_lut_3_lut (.I0(\Gain1_mul_temp[4] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[4] ), .I3(GND_net), 
            .O(n9));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i9_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i5_3_lut_4_lut (.I0(\Gain1_mul_temp[4] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[4] ), .O(\Max_out1[4] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i5_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 in0_2_31__I_0_i4_3_lut_4_lut (.I0(\Gain1_mul_temp[3] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(out0_31__N_334), .I3(\abcVoltage_2[3] ), .O(\Max_out1[3] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_2_31__I_0_i4_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 Max_stage1_val_0__31__I_0_i7_2_lut_3_lut (.I0(\Gain1_mul_temp[3] ), 
            .I1(Max_stage1_val_0__31__N_335), .I2(\abcVoltage_2[3] ), .I3(GND_net), 
            .O(n7));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam Max_stage1_val_0__31__I_0_i7_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 in0_2_31__I_0_i16_3_lut (.I0(\abcVoltage_2[15] ), .I1(\Max_stage1_val[0] [15]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[15] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i17_3_lut (.I0(\abcVoltage_2[16] ), .I1(\Max_stage1_val[0] [16]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[16] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i18_3_lut (.I0(\abcVoltage_2[17] ), .I1(\Max_stage1_val[0] [17]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[17] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i19_3_lut (.I0(\abcVoltage_2[18] ), .I1(\Max_stage1_val[0] [18]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[18] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i32_3_lut (.I0(\abcVoltage_2[31] ), .I1(\Max_stage1_val[0] [31]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[31] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i20_3_lut (.I0(\abcVoltage_2[19] ), .I1(\Max_stage1_val[0] [19]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[19] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i21_3_lut (.I0(\abcVoltage_2[20] ), .I1(\Max_stage1_val[0] [20]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[20] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i22_3_lut (.I0(\abcVoltage_2[21] ), .I1(\Max_stage1_val[0] [21]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[21] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i23_3_lut (.I0(\abcVoltage_2[22] ), .I1(\Max_stage1_val[0] [22]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[22] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i24_3_lut (.I0(\abcVoltage_2[23] ), .I1(\Max_stage1_val[0] [23]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[23] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i25_3_lut (.I0(\abcVoltage_2[24] ), .I1(\Max_stage1_val[0] [24]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[24] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i26_3_lut (.I0(\abcVoltage_2[25] ), .I1(\Max_stage1_val[0] [25]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[25] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i27_3_lut (.I0(\abcVoltage_2[26] ), .I1(\Max_stage1_val[0] [26]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[26] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i28_3_lut (.I0(\abcVoltage_2[27] ), .I1(\Max_stage1_val[0] [27]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[27] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i29_3_lut (.I0(\abcVoltage_2[28] ), .I1(\Max_stage1_val[0] [28]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[28] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i30_3_lut (.I0(\abcVoltage_2[29] ), .I1(\Max_stage1_val[0] [29]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[29] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_2_31__I_0_i31_3_lut (.I0(\abcVoltage_2[30] ), .I1(\Max_stage1_val[0] [30]), 
            .I2(out0_31__N_334), .I3(GND_net), .O(\Max_out1[30] ));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[27] 53[33])
    defparam in0_2_31__I_0_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i30_3_lut (.I0(\abcVoltage_1[29] ), .I1(alphaVoltage[14]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [29]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i31_3_lut (.I0(\abcVoltage_1[30] ), .I1(alphaVoltage[15]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [30]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i29_3_lut (.I0(\abcVoltage_1[28] ), .I1(alphaVoltage[13]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [28]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i28_3_lut (.I0(\abcVoltage_1[27] ), .I1(alphaVoltage[12]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [27]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i27_3_lut (.I0(\abcVoltage_1[26] ), .I1(alphaVoltage[11]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [26]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i24_rep_81_3_lut (.I0(\abcVoltage_1[23] ), .I1(alphaVoltage[8]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [23]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i24_rep_81_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i47_2_lut (.I0(\abcVoltage_2[23] ), 
            .I1(\Max_stage1_val[0] [23]), .I2(GND_net), .I3(GND_net), 
            .O(n47));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i47_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Max_stage1_val_0__31__I_0_i45_2_lut (.I0(\abcVoltage_2[22] ), 
            .I1(\Max_stage1_val[0] [22]), .I2(GND_net), .I3(GND_net), 
            .O(n45));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i23_rep_80_3_lut (.I0(\abcVoltage_1[22] ), .I1(alphaVoltage[7]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [22]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i23_rep_80_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i19_rep_76_3_lut (.I0(\abcVoltage_1[18] ), .I1(alphaVoltage[3]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [18]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i19_rep_76_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i18_rep_75_3_lut (.I0(\abcVoltage_1[17] ), .I1(alphaVoltage[2]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [17]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i18_rep_75_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i17_rep_74_3_lut (.I0(\abcVoltage_1[16] ), .I1(alphaVoltage[1]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [16]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i17_rep_74_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i33_2_lut (.I0(\abcVoltage_2[16] ), 
            .I1(\Max_stage1_val[0] [16]), .I2(GND_net), .I3(GND_net), 
            .O(n33));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Max_stage1_val_0__31__I_0_i35_2_lut (.I0(\abcVoltage_2[17] ), 
            .I1(\Max_stage1_val[0] [17]), .I2(GND_net), .I3(GND_net), 
            .O(n35));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Max_stage1_val_0__31__I_0_i37_2_lut (.I0(\abcVoltage_2[18] ), 
            .I1(\Max_stage1_val[0] [18]), .I2(GND_net), .I3(GND_net), 
            .O(n37));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i16_rep_73_3_lut (.I0(\abcVoltage_1[15] ), .I1(alphaVoltage[0]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [15]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i16_rep_73_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i31_2_lut (.I0(\abcVoltage_2[15] ), 
            .I1(\Max_stage1_val[0] [15]), .I2(GND_net), .I3(GND_net), 
            .O(n31));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13110_2_lut (.I0(\Gain1_mul_temp[1] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(GND_net), .I3(GND_net), .O(\Max_stage1_val[0] [1]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam i13110_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13111_2_lut (.I0(\Gain1_mul_temp[2] ), .I1(Max_stage1_val_0__31__N_335), 
            .I2(GND_net), .I3(GND_net), .O(\Max_stage1_val[0] [2]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam i13111_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 in0_0_31__I_0_i40_3_lut (.I0(n38), .I1(alphaVoltage[6]), .I2(n43), 
            .I3(GND_net), .O(n40));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16900_3_lut (.I0(n56), .I1(n40), .I2(n21842), .I3(GND_net), 
            .O(n21912));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16902_3_lut (.I0(n52), .I1(n21912), .I2(n21844), .I3(GND_net), 
            .O(n21914));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i22_rep_79_3_lut (.I0(\abcVoltage_1[21] ), .I1(alphaVoltage[6]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [21]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i22_rep_79_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i21_rep_78_3_lut (.I0(\abcVoltage_1[20] ), .I1(alphaVoltage[5]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [20]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i21_rep_78_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_1_31__I_0_i20_rep_77_3_lut (.I0(\abcVoltage_1[19] ), .I1(alphaVoltage[4]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [19]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i20_rep_77_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i39_2_lut (.I0(\abcVoltage_2[19] ), 
            .I1(\Max_stage1_val[0] [19]), .I2(GND_net), .I3(GND_net), 
            .O(n39));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Max_stage1_val_0__31__I_0_i41_2_lut (.I0(\abcVoltage_2[20] ), 
            .I1(\Max_stage1_val[0] [20]), .I2(GND_net), .I3(GND_net), 
            .O(n41));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Max_stage1_val_0__31__I_0_i43_2_lut (.I0(\abcVoltage_2[21] ), 
            .I1(\Max_stage1_val[0] [21]), .I2(GND_net), .I3(GND_net), 
            .O(n43_adj_2183));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i26_3_lut (.I0(\abcVoltage_1[25] ), .I1(alphaVoltage[10]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [25]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i51_2_lut (.I0(\abcVoltage_2[25] ), 
            .I1(\Max_stage1_val[0] [25]), .I2(GND_net), .I3(GND_net), 
            .O(n51));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i51_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Max_stage1_val_0__31__I_0_i49_2_lut (.I0(\abcVoltage_2[24] ), 
            .I1(\Max_stage1_val[0] [24]), .I2(GND_net), .I3(GND_net), 
            .O(n49));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i49_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_1_31__I_0_i25_3_lut (.I0(\abcVoltage_1[24] ), .I1(alphaVoltage[9]), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(\Max_stage1_val[0] [24]));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[30] 46[22])
    defparam in0_1_31__I_0_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_0_31__I_0_i49_2_lut (.I0(\abcVoltage_1[24] ), .I1(alphaVoltage[9]), 
            .I2(GND_net), .I3(GND_net), .O(n49_adj_2184));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i49_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i51_2_lut (.I0(\abcVoltage_1[25] ), .I1(alphaVoltage[10]), 
            .I2(GND_net), .I3(GND_net), .O(n51_adj_2185));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i51_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i53_2_lut (.I0(\abcVoltage_1[26] ), .I1(alphaVoltage[11]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i53_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i45_2_lut (.I0(\abcVoltage_1[22] ), .I1(alphaVoltage[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_2186));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i47_2_lut (.I0(\abcVoltage_1[23] ), .I1(alphaVoltage[8]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_2187));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i47_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i37_2_lut (.I0(\abcVoltage_1[18] ), .I1(alphaVoltage[3]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_2188));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16718_4_lut (.I0(n41_adj_2189), .I1(n39_adj_2190), .I2(n37_adj_2188), 
            .I3(n21545), .O(n21730));
    defparam i16718_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i16537_4_lut (.I0(n47_adj_2187), .I1(n45_adj_2186), .I2(n43), 
            .I3(n21730), .O(n21549));
    defparam i16537_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i16914_4_lut (.I0(n53), .I1(n51_adj_2185), .I2(n49_adj_2184), 
            .I3(n21549), .O(n21926));
    defparam i16914_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16832_4_lut (.I0(n59), .I1(n57), .I2(n55), .I3(n21926), 
            .O(n21844));
    defparam i16832_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 in0_0_31__I_0_i36_3_lut (.I0(alphaVoltage[3]), .I1(alphaVoltage[7]), 
            .I2(n45_adj_2186), .I3(GND_net), .O(n36));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_0_31__I_0_i44_3_lut (.I0(n36), .I1(alphaVoltage[8]), .I2(n47_adj_2187), 
            .I3(GND_net), .O(n44));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i44_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16997_4_lut (.I0(n44), .I1(n34), .I2(n47_adj_2187), .I3(n21547), 
            .O(n22009));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16997_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i16998_3_lut (.I0(n22009), .I1(alphaVoltage[9]), .I2(n49_adj_2184), 
            .I3(GND_net), .O(n22010));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16949_3_lut (.I0(n22010), .I1(alphaVoltage[10]), .I2(n51_adj_2185), 
            .I3(GND_net), .O(n21961));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16663_3_lut (.I0(n21961), .I1(alphaVoltage[11]), .I2(n53), 
            .I3(GND_net), .O(n52));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_0_31__I_0_i55_2_lut (.I0(\abcVoltage_1[27] ), .I1(alphaVoltage[12]), 
            .I2(GND_net), .I3(GND_net), .O(n55));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i55_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i57_2_lut (.I0(\abcVoltage_1[28] ), .I1(alphaVoltage[13]), 
            .I2(GND_net), .I3(GND_net), .O(n57));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i57_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i59_2_lut (.I0(\abcVoltage_1[29] ), .I1(alphaVoltage[14]), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i59_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i39_2_lut (.I0(\abcVoltage_1[19] ), .I1(alphaVoltage[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_2190));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i41_2_lut (.I0(\abcVoltage_1[20] ), .I1(alphaVoltage[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_2189));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16648_3_lut (.I0(n43), .I1(n41_adj_2189), .I2(n39_adj_2190), 
            .I3(GND_net), .O(n21660));
    defparam i16648_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i16830_4_lut (.I0(n59), .I1(n57), .I2(n55), .I3(n21660), 
            .O(n21842));
    defparam i16830_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut (.I0(\Gain1_mul_temp[4] ), .I1(\Gain1_mul_temp[3] ), 
            .I2(\Gain1_mul_temp[2] ), .I3(\Gain1_mul_temp[1] ), .O(n20038));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_309 (.I0(\Gain1_mul_temp[7] ), .I1(\Gain1_mul_temp[6] ), 
            .I2(\Gain1_mul_temp[5] ), .I3(n20038), .O(n20044));
    defparam i1_4_lut_adj_309.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_310 (.I0(\Gain1_mul_temp[10] ), .I1(\Gain1_mul_temp[9] ), 
            .I2(\Gain1_mul_temp[8] ), .I3(n20044), .O(n20050));
    defparam i1_4_lut_adj_310.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_311 (.I0(\Gain1_mul_temp[13] ), .I1(\Gain1_mul_temp[12] ), 
            .I2(\Gain1_mul_temp[11] ), .I3(n20050), .O(n20056));
    defparam i1_4_lut_adj_311.LUT_INIT = 16'hfffe;
    SB_LUT4 in0_0_31__I_0_i32_4_lut (.I0(n20056), .I1(alphaVoltage[0]), 
            .I2(\abcVoltage_1[15] ), .I3(\abcVoltage_1[14] ), .O(n32));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i32_4_lut.LUT_INIT = 16'h0c4d;
    SB_LUT4 i16868_3_lut (.I0(n32), .I1(alphaVoltage[12]), .I2(n55), .I3(GND_net), 
            .O(n21880));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16869_3_lut (.I0(n21880), .I1(alphaVoltage[13]), .I2(n57), 
            .I3(GND_net), .O(n21881));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16665_3_lut (.I0(n21881), .I1(alphaVoltage[14]), .I2(n59), 
            .I3(GND_net), .O(n56));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam i16665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 in0_0_31__I_0_i43_2_lut (.I0(\abcVoltage_1[21] ), .I1(alphaVoltage[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 in0_0_31__I_0_i38_3_lut (.I0(alphaVoltage[4]), .I1(alphaVoltage[5]), 
            .I2(n41_adj_2189), .I3(GND_net), .O(n38));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(45[31:47])
    defparam in0_0_31__I_0_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16635_3_lut (.I0(n27), .I1(n25), .I2(n23), .I3(GND_net), 
            .O(n21647));
    defparam i16635_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 Max_stage1_val_0__31__I_0_i20_3_lut (.I0(\Gain1_mul_temp[11] ), 
            .I1(\Gain1_mul_temp[12] ), .I2(n25), .I3(GND_net), .O(n21515));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16756_3_lut (.I0(n51), .I1(n49), .I2(n27), .I3(GND_net), 
            .O(n21768));
    defparam i16756_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 Max_stage1_val_0__31__I_0_i44_3_lut (.I0(n22), .I1(\Max_stage1_val[0] [25]), 
            .I2(n51), .I3(GND_net), .O(n44_adj_2191));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i44_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16768_3_lut (.I0(n21), .I1(n19), .I2(n11), .I3(GND_net), 
            .O(n21780));
    defparam i16768_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i16812_4_lut (.I0(n27), .I1(n25), .I2(n23), .I3(n21780), 
            .O(n21824));
    defparam i16812_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i16870_4_lut (.I0(n43_adj_2183), .I1(n41), .I2(n39), .I3(n21824), 
            .O(n21882));
    defparam i16870_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i16626_4_lut (.I0(n29), .I1(n17), .I2(n15), .I3(n13), .O(n21638));
    defparam i16626_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i4_5_3_lut (.I0(\abcVoltage_2[1] ), .I1(\Gain1_mul_temp[1] ), 
            .I2(Max_stage1_val_0__31__N_335), .I3(GND_net), .O(n19887));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i4_5_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 Max_stage1_val_0__31__I_0_i6_4_lut (.I0(n19887), .I1(\Max_stage1_val[0] [2]), 
            .I2(\abcVoltage_2[2] ), .I3(\Max_stage1_val[0] [1]), .O(n6));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i6_4_lut.LUT_INIT = 16'hcf4d;
    SB_LUT4 i16491_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n7), .O(n21497));
    defparam i16491_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16620_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n21497), 
            .O(n21632));
    defparam i16620_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16926_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n21632), 
            .O(n21938));
    defparam i16926_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16808_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n21938), 
            .O(n21820));
    defparam i16808_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i17001_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n21820), 
            .O(n22013));
    defparam i17001_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16878_4_lut (.I0(n43_adj_2183), .I1(n41), .I2(n39), .I3(n22013), 
            .O(n21890));
    defparam i16878_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 Max_stage1_val_0__31__I_0_i10_3_lut (.I0(\Gain1_mul_temp[5] ), 
            .I1(\Gain1_mul_temp[9] ), .I2(n19), .I3(GND_net), .O(n21507));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i18_3_lut (.I0(n21507), .I1(\Gain1_mul_temp[10] ), 
            .I2(n21), .I3(GND_net), .O(n21513));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i8_3_lut (.I0(\Gain1_mul_temp[3] ), 
            .I1(\Gain1_mul_temp[4] ), .I2(n9), .I3(GND_net), .O(n21505));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16575_4_lut (.I0(n49), .I1(n47), .I2(n45), .I3(n21647), 
            .O(n21587));
    defparam i16575_4_lut.LUT_INIT = 16'habaa;
    SB_LUT4 i16975_4_lut (.I0(n44_adj_2191), .I1(Max_stage1_val_0__31__N_335), 
            .I2(n21768), .I3(n21515), .O(n21987));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16975_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 Max_stage1_val_0__31__I_0_i42_3_lut (.I0(n24), .I1(\Max_stage1_val[0] [23]), 
            .I2(n47), .I3(GND_net), .O(n42));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16945_3_lut (.I0(n21956), .I1(\Max_stage1_val[0] [20]), .I2(n41), 
            .I3(GND_net), .O(n21957));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16856_4_lut (.I0(n49), .I1(n47), .I2(n45), .I3(n21882), 
            .O(n21868));
    defparam i16856_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i17029_4_lut (.I0(n42), .I1(n21987), .I2(n51), .I3(n21587), 
            .O(n22041));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17029_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16669_3_lut (.I0(n21957), .I1(\Max_stage1_val[0] [21]), .I2(n43_adj_2183), 
            .I3(GND_net), .O(n21681));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i12_3_lut (.I0(\Gain1_mul_temp[6] ), 
            .I1(\Gain1_mul_temp[7] ), .I2(n15), .I3(GND_net), .O(n21509));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Max_stage1_val_0__31__I_0_i14_3_lut (.I0(n21509), .I1(\Gain1_mul_temp[8] ), 
            .I2(n17), .I3(GND_net), .O(n21511));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16947_3_lut (.I0(n21958), .I1(\Max_stage1_val[0] [17]), .I2(n35), 
            .I3(GND_net), .O(n21959));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16802_4_lut (.I0(n35), .I1(n33), .I2(n31), .I3(n21638), 
            .O(n21814));
    defparam i16802_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i17027_3_lut (.I0(n16), .I1(\Max_stage1_val[0] [15]), .I2(n31), 
            .I3(GND_net), .O(n22039));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16667_3_lut (.I0(n21959), .I1(\Max_stage1_val[0] [18]), .I2(n37), 
            .I3(GND_net), .O(n21679));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17025_4_lut (.I0(n49), .I1(n47), .I2(n45), .I3(n21890), 
            .O(n22037));
    defparam i17025_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17060_4_lut (.I0(n21681), .I1(n22041), .I2(n51), .I3(n21868), 
            .O(n22072));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17060_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i17048_4_lut (.I0(n21679), .I1(n22039), .I2(n37), .I3(n21814), 
            .O(n22060));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17048_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i17075_4_lut (.I0(n22060), .I1(n22072), .I2(n51), .I3(n22037), 
            .O(n22087));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17075_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i17076_3_lut (.I0(n22087), .I1(\Max_stage1_val[0] [26]), .I2(\abcVoltage_2[26] ), 
            .I3(GND_net), .O(n22088));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17076_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i17074_3_lut (.I0(n22088), .I1(\Max_stage1_val[0] [27]), .I2(\abcVoltage_2[27] ), 
            .I3(GND_net), .O(n22086));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17074_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i17062_3_lut (.I0(n22086), .I1(\Max_stage1_val[0] [28]), .I2(\abcVoltage_2[28] ), 
            .I3(GND_net), .O(n22074));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17062_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i17063_3_lut (.I0(n22074), .I1(\Max_stage1_val[0] [29]), .I2(\abcVoltage_2[29] ), 
            .I3(GND_net), .O(n22075));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17063_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i17051_3_lut (.I0(n22075), .I1(\Max_stage1_val[0] [30]), .I2(\abcVoltage_2[30] ), 
            .I3(GND_net), .O(n22063));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17051_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i17012_3_lut (.I0(n22063), .I1(\abcVoltage_2[31] ), .I2(\Max_stage1_val[0] [31]), 
            .I3(GND_net), .O(out0_31__N_334));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i17012_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16946_4_lut_4_lut (.I0(Max_stage1_val_0__31__N_335), .I1(\Max_stage1_val[0] [16]), 
            .I2(\abcVoltage_2[16] ), .I3(n21511), .O(n21958));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16946_4_lut_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 Max_stage1_val_0__31__I_0_i24_4_lut_4_lut (.I0(Max_stage1_val_0__31__N_335), 
            .I1(\Max_stage1_val[0] [22]), .I2(\abcVoltage_2[22] ), .I3(n21505), 
            .O(n24));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam Max_stage1_val_0__31__I_0_i24_4_lut_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i16944_4_lut_4_lut (.I0(Max_stage1_val_0__31__N_335), .I1(\Max_stage1_val[0] [19]), 
            .I2(\abcVoltage_2[19] ), .I3(n21513), .O(n21956));   // ../../hdlcoderFocCurrentFixptHdl/Max.v(52[28:66])
    defparam i16944_4_lut_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i16535_2_lut_4_lut (.I0(\abcVoltage_1[22] ), .I1(alphaVoltage[7]), 
            .I2(\abcVoltage_1[18] ), .I3(alphaVoltage[3]), .O(n21547));
    defparam i16535_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    
endmodule
//
// Verilog Description of module Sine_Cosine
//

module Sine_Cosine (GND_net, \Amp25_out1[14] , \Product_mul_temp[26] , 
            Look_Up_Table_out1_1) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \Amp25_out1[14] ;
    input \Product_mul_temp[26] ;
    output [15:0]Look_Up_Table_out1_1;
    
    
    Sine_Cosine_LUT u_Sine_Cosine_LUT (.GND_net(GND_net), .\Amp25_out1[14] (\Amp25_out1[14] ), 
            .\Product_mul_temp[26] (\Product_mul_temp[26] ), .Look_Up_Table_out1_1({Look_Up_Table_out1_1})) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine.v(43[19] 46[39])
    
endmodule
//
// Verilog Description of module Sine_Cosine_LUT
//

module Sine_Cosine_LUT (GND_net, \Amp25_out1[14] , \Product_mul_temp[26] , 
            Look_Up_Table_out1_1) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \Amp25_out1[14] ;
    input \Product_mul_temp[26] ;
    output [15:0]Look_Up_Table_out1_1;
    
    wire [31:0]n3374;
    wire [31:0]n3375;
    
    wire n17429, n17423, n2828, n17424, n17422, n17421;
    wire [15:0]Look_Up_Table_sub_temp1;   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(103[21:44])
    
    wire n17432;
    wire [31:0]n3376;
    
    wire n2831, n17433;
    wire [31:0]n3373;
    
    wire n17419, n3236, n2825, n17418, n17417, n17416, n17415, 
        n17414, n17413, n17412, n15467, n15468, n15469, n2834, 
        n15470, n2840, n15466, VCC_net, n15471, n2843, n2810, 
        n15460, n2807;
    wire [31:0]n3372;
    
    wire n17410, n3232, n2822, n17409, n17408, n17407, n17406, 
        n17405, n17404, n17403;
    wire [31:0]n3371;
    
    wire n17401, n3228, n2819, n17400, n17399, n15465, n17398, 
        n15461, n17397, n15464, n17396, n17395, n17394;
    wire [31:0]n3370;
    
    wire n17392, n3224, n2816, n17391, n17390, n17389, n17388, 
        n17387, n17386, n17385;
    wire [31:0]n3369;
    
    wire n17383, n3220, n2813, n17382, n17381, n17380, n17379, 
        n17378, n17377, n17376;
    wire [31:0]n3368;
    
    wire n17374, n3216, n17373, n17372, n17371, n17370, n17369, 
        n17368, n17367;
    wire [31:0]n3367;
    
    wire n17365, n3212, n17364, n17363, n17362, n17361, n17360, 
        n17359, n17358;
    wire [8:0]n7464;
    wire [7:0]n7546;
    
    wire n2652, n17357, n17356, n17355, n17354, n17353, n17352, 
        n17351, n15463, n17350;
    wire [6:0]n7890;
    wire [5:0]n8171;
    
    wire n17349, n17348, n17431, n17347, n17346, n17345, n17344, 
        n17343, n17342, n17341, n17340, n17339, n17338, n17337;
    wire [4:0]n8488;
    
    wire n17336, n17335, n17334, n17333, n17332, n3240, n17428, 
        n15462;
    wire [48:0]Look_Up_Table_mul_temp1;   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(104[21:44])
    wire [31:0]n3380;
    
    wire n3260, n17504;
    wire [31:0]n3379;
    
    wire n3256, n17503;
    wire [31:0]n3378;
    
    wire n3252, n17502;
    wire [31:0]n3377;
    
    wire n3248, n17501, n3244, n17500, n17499, n17498, n17497, 
        n17496, n17495, n17494, n17493, n17492, n17491, n17490, 
        n17489, n17488, n17487, n17486, n17485, n17484, n17483, 
        n17482, n17481, n17479, n17478, n17477, n17476, n17475, 
        n17474, n17473, n17472, n17471, n17469, n17468, n17467, 
        n17466, n17465, n17464, n17463, n17462, n17461, n17459, 
        n17458, n17457, n17456, n17455, n17454, n17453, n17452, 
        n17451, n17449, n17448, n17447, n17446, n17445, n17444, 
        n17443, n17442, n17441, n17439, n17427, n17426, n17425, 
        n17438, n17437, n15956, n15955, n15954, n15953, n15952, 
        n15951, n15950, n15949, n15948, n15947, n15946, n15945, 
        n15944, n17436, n17435, n17434;
    
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_11_lut (.I0(GND_net), .I1(n3375[30]), 
            .I2(GND_net), .I3(n17429), .O(n3374[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_5 (.CI(n17423), .I0(n3375[24]), 
            .I1(n2828), .CO(n17424));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_4_lut (.I0(GND_net), .I1(n3375[23]), 
            .I2(n2828), .I3(n17422), .O(n3374[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_4 (.CI(n17422), .I0(n3375[23]), 
            .I1(n2828), .CO(n17423));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_3_lut (.I0(GND_net), .I1(n3375[22]), 
            .I2(GND_net), .I3(n17421), .O(n3374[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_3 (.CI(n17421), .I0(n3375[22]), 
            .I1(GND_net), .CO(n17422));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2828), .I3(GND_net), .O(n3374[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2828), .CO(n17421));
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_4 (.CI(n17432), .I0(n3376[23]), 
            .I1(n2831), .CO(n17433));
    SB_LUT4 add_5961_10_lut (.I0(GND_net), .I1(n3374[30]), .I2(GND_net), 
            .I3(n17419), .O(n3373[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_10 (.CI(n17419), .I0(n3374[30]), .I1(GND_net), .CO(n3236));
    SB_LUT4 add_5961_9_lut (.I0(GND_net), .I1(n3374[29]), .I2(n2825), 
            .I3(n17418), .O(n3373[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_9 (.CI(n17418), .I0(n3374[29]), .I1(n2825), .CO(n17419));
    SB_LUT4 add_5961_8_lut (.I0(GND_net), .I1(n3374[28]), .I2(n2825), 
            .I3(n17417), .O(n3373[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_8 (.CI(n17417), .I0(n3374[28]), .I1(n2825), .CO(n17418));
    SB_LUT4 add_5961_7_lut (.I0(GND_net), .I1(n3374[27]), .I2(n2825), 
            .I3(n17416), .O(n3373[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_7 (.CI(n17416), .I0(n3374[27]), .I1(n2825), .CO(n17417));
    SB_LUT4 add_5961_6_lut (.I0(GND_net), .I1(n3374[26]), .I2(n2825), 
            .I3(n17415), .O(n3373[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_6 (.CI(n17415), .I0(n3374[26]), .I1(n2825), .CO(n17416));
    SB_LUT4 add_5961_5_lut (.I0(GND_net), .I1(n3374[25]), .I2(n2825), 
            .I3(n17414), .O(n3373[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_5 (.CI(n17414), .I0(n3374[25]), .I1(n2825), .CO(n17415));
    SB_LUT4 add_5961_4_lut (.I0(GND_net), .I1(n3374[24]), .I2(n2825), 
            .I3(n17413), .O(n3373[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_4 (.CI(n17413), .I0(n3374[24]), .I1(n2825), .CO(n17414));
    SB_LUT4 add_5961_3_lut (.I0(GND_net), .I1(n3374[23]), .I2(n2825), 
            .I3(n17412), .O(n3373[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_10 (.CI(n15467), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15468));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15467), .O(n2831)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_11 (.CI(n15468), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15469));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15468), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_12 (.CI(n15469), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15470));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15469), .O(n2840)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15466), .O(n2828)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_13 (.CI(n15470), .I0(VCC_net), 
            .I1(\Product_mul_temp[26] ), .CO(n15471));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut (.I0(\Product_mul_temp[26] ), 
            .I1(VCC_net), .I2(\Product_mul_temp[26] ), .I3(n15470), .O(n2843)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_9 (.CI(n15466), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15467));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(VCC_net), .I3(n15471), .O(Look_Up_Table_sub_temp1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_3 (.CI(n17412), .I0(n3374[23]), .I1(n2825), .CO(n17413));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15460), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(VCC_net), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_5961_2_lut (.I0(GND_net), .I1(n3374[22]), .I2(GND_net), 
            .I3(GND_net), .O(n3373[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5961_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5961_2 (.CI(GND_net), .I0(n3374[22]), .I1(GND_net), .CO(n17412));
    SB_LUT4 add_5960_10_lut (.I0(GND_net), .I1(n3373[30]), .I2(GND_net), 
            .I3(n17410), .O(n3372[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_10 (.CI(n17410), .I0(n3373[30]), .I1(GND_net), .CO(n3232));
    SB_LUT4 add_5960_9_lut (.I0(GND_net), .I1(n3373[29]), .I2(n2822), 
            .I3(n17409), .O(n3372[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_9 (.CI(n17409), .I0(n3373[29]), .I1(n2822), .CO(n17410));
    SB_LUT4 add_5960_8_lut (.I0(GND_net), .I1(n3373[28]), .I2(n2822), 
            .I3(n17408), .O(n3372[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_8 (.CI(n17408), .I0(n3373[28]), .I1(n2822), .CO(n17409));
    SB_LUT4 add_5960_7_lut (.I0(GND_net), .I1(n3373[27]), .I2(n2822), 
            .I3(n17407), .O(n3372[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_7 (.CI(n17407), .I0(n3373[27]), .I1(n2822), .CO(n17408));
    SB_LUT4 add_5960_6_lut (.I0(GND_net), .I1(n3373[26]), .I2(n2822), 
            .I3(n17406), .O(n3372[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_6 (.CI(n17406), .I0(n3373[26]), .I1(n2822), .CO(n17407));
    SB_LUT4 add_5960_5_lut (.I0(GND_net), .I1(n3373[25]), .I2(n2822), 
            .I3(n17405), .O(n3372[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_5 (.CI(n17405), .I0(n3373[25]), .I1(n2822), .CO(n17406));
    SB_LUT4 add_5960_4_lut (.I0(GND_net), .I1(n3373[24]), .I2(n2822), 
            .I3(n17404), .O(n3372[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_4 (.CI(n17404), .I0(n3373[24]), .I1(n2822), .CO(n17405));
    SB_LUT4 add_5960_3_lut (.I0(GND_net), .I1(n3373[23]), .I2(n2822), 
            .I3(n17403), .O(n3372[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_3 (.CI(n17403), .I0(n3373[23]), .I1(n2822), .CO(n17404));
    SB_LUT4 add_5960_2_lut (.I0(GND_net), .I1(n2825), .I2(GND_net), .I3(GND_net), 
            .O(n3372[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5960_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5960_2 (.CI(GND_net), .I0(n2825), .I1(GND_net), .CO(n17403));
    SB_LUT4 add_5959_10_lut (.I0(GND_net), .I1(n3372[30]), .I2(GND_net), 
            .I3(n17401), .O(n3371[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_10 (.CI(n17401), .I0(n3372[30]), .I1(GND_net), .CO(n3228));
    SB_LUT4 add_5959_9_lut (.I0(GND_net), .I1(n3372[29]), .I2(n2819), 
            .I3(n17400), .O(n3371[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_9 (.CI(n17400), .I0(n3372[29]), .I1(n2819), .CO(n17401));
    SB_LUT4 add_5959_8_lut (.I0(GND_net), .I1(n3372[28]), .I2(n2819), 
            .I3(n17399), .O(n3371[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15465), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15460));
    SB_CARRY add_5959_8 (.CI(n17399), .I0(n3372[28]), .I1(n2819), .CO(n17400));
    SB_LUT4 add_5959_7_lut (.I0(GND_net), .I1(n3372[27]), .I2(n2819), 
            .I3(n17398), .O(n3371[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_7 (.CI(n17398), .I0(n3372[27]), .I1(n2819), .CO(n17399));
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_3 (.CI(n15460), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15461));
    SB_LUT4 add_5959_6_lut (.I0(GND_net), .I1(n3372[26]), .I2(n2819), 
            .I3(n17397), .O(n3371[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_8 (.CI(n15465), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15466));
    SB_CARRY add_5959_6 (.CI(n17397), .I0(n3372[26]), .I1(n2819), .CO(n17398));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15464), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_5959_5_lut (.I0(GND_net), .I1(n3372[25]), .I2(n2819), 
            .I3(n17396), .O(n3371[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_5 (.CI(n17396), .I0(n3372[25]), .I1(n2819), .CO(n17397));
    SB_LUT4 add_5959_4_lut (.I0(GND_net), .I1(n3372[24]), .I2(n2819), 
            .I3(n17395), .O(n3371[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_4 (.CI(n17395), .I0(n3372[24]), .I1(n2819), .CO(n17396));
    SB_LUT4 add_5959_3_lut (.I0(GND_net), .I1(n3372[23]), .I2(n2819), 
            .I3(n17394), .O(n3371[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_3 (.CI(n17394), .I0(n3372[23]), .I1(n2819), .CO(n17395));
    SB_LUT4 add_5959_2_lut (.I0(GND_net), .I1(n2822), .I2(GND_net), .I3(GND_net), 
            .O(n3371[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5959_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5959_2 (.CI(GND_net), .I0(n2822), .I1(GND_net), .CO(n17394));
    SB_LUT4 add_5958_10_lut (.I0(GND_net), .I1(n3371[30]), .I2(GND_net), 
            .I3(n17392), .O(n3370[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_10 (.CI(n17392), .I0(n3371[30]), .I1(GND_net), .CO(n3224));
    SB_LUT4 add_5958_9_lut (.I0(GND_net), .I1(n3371[29]), .I2(n2816), 
            .I3(n17391), .O(n3370[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_9 (.CI(n17391), .I0(n3371[29]), .I1(n2816), .CO(n17392));
    SB_LUT4 add_5958_8_lut (.I0(GND_net), .I1(n3371[28]), .I2(n2816), 
            .I3(n17390), .O(n3370[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_8 (.CI(n17390), .I0(n3371[28]), .I1(n2816), .CO(n17391));
    SB_LUT4 add_5958_7_lut (.I0(GND_net), .I1(n3371[27]), .I2(n2816), 
            .I3(n17389), .O(n3370[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_7 (.CI(n17389), .I0(n3371[27]), .I1(n2816), .CO(n17390));
    SB_LUT4 add_5958_6_lut (.I0(GND_net), .I1(n3371[26]), .I2(n2816), 
            .I3(n17388), .O(n3370[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_6 (.CI(n17388), .I0(n3371[26]), .I1(n2816), .CO(n17389));
    SB_LUT4 add_5958_5_lut (.I0(GND_net), .I1(n3371[25]), .I2(n2816), 
            .I3(n17387), .O(n3370[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_5 (.CI(n17387), .I0(n3371[25]), .I1(n2816), .CO(n17388));
    SB_LUT4 add_5958_4_lut (.I0(GND_net), .I1(n3371[24]), .I2(n2816), 
            .I3(n17386), .O(n3370[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_4 (.CI(n17386), .I0(n3371[24]), .I1(n2816), .CO(n17387));
    SB_LUT4 add_5958_3_lut (.I0(GND_net), .I1(n3371[23]), .I2(n2816), 
            .I3(n17385), .O(n3370[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_3 (.CI(n17385), .I0(n3371[23]), .I1(n2816), .CO(n17386));
    SB_LUT4 add_5958_2_lut (.I0(GND_net), .I1(n2819), .I2(GND_net), .I3(GND_net), 
            .O(n3370[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5958_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5958_2 (.CI(GND_net), .I0(n2819), .I1(GND_net), .CO(n17385));
    SB_LUT4 add_5957_10_lut (.I0(GND_net), .I1(n3370[30]), .I2(GND_net), 
            .I3(n17383), .O(n3369[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_10 (.CI(n17383), .I0(n3370[30]), .I1(GND_net), .CO(n3220));
    SB_LUT4 add_5957_9_lut (.I0(GND_net), .I1(n3370[29]), .I2(n2813), 
            .I3(n17382), .O(n3369[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_9 (.CI(n17382), .I0(n3370[29]), .I1(n2813), .CO(n17383));
    SB_LUT4 add_5957_8_lut (.I0(GND_net), .I1(n3370[28]), .I2(n2813), 
            .I3(n17381), .O(n3369[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_8 (.CI(n17381), .I0(n3370[28]), .I1(n2813), .CO(n17382));
    SB_LUT4 add_5957_7_lut (.I0(GND_net), .I1(n3370[27]), .I2(n2813), 
            .I3(n17380), .O(n3369[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_7 (.CI(n17380), .I0(n3370[27]), .I1(n2813), .CO(n17381));
    SB_LUT4 add_5957_6_lut (.I0(GND_net), .I1(n3370[26]), .I2(n2813), 
            .I3(n17379), .O(n3369[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_6 (.CI(n17379), .I0(n3370[26]), .I1(n2813), .CO(n17380));
    SB_LUT4 add_5957_5_lut (.I0(GND_net), .I1(n3370[25]), .I2(n2813), 
            .I3(n17378), .O(n3369[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_5 (.CI(n17378), .I0(n3370[25]), .I1(n2813), .CO(n17379));
    SB_LUT4 add_5957_4_lut (.I0(GND_net), .I1(n3370[24]), .I2(n2813), 
            .I3(n17377), .O(n3369[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_4 (.CI(n17377), .I0(n3370[24]), .I1(n2813), .CO(n17378));
    SB_LUT4 add_5957_3_lut (.I0(GND_net), .I1(n3370[23]), .I2(n2813), 
            .I3(n17376), .O(n3369[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_3 (.CI(n17376), .I0(n3370[23]), .I1(n2813), .CO(n17377));
    SB_LUT4 add_5957_2_lut (.I0(GND_net), .I1(n2816), .I2(GND_net), .I3(GND_net), 
            .O(n3369[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_2 (.CI(GND_net), .I0(n2816), .I1(GND_net), .CO(n17376));
    SB_LUT4 add_5956_10_lut (.I0(GND_net), .I1(n3369[30]), .I2(GND_net), 
            .I3(n17374), .O(n3368[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_10 (.CI(n17374), .I0(n3369[30]), .I1(GND_net), .CO(n3216));
    SB_LUT4 add_5956_9_lut (.I0(GND_net), .I1(n3369[29]), .I2(n2810), 
            .I3(n17373), .O(n3368[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_9 (.CI(n17373), .I0(n3369[29]), .I1(n2810), .CO(n17374));
    SB_LUT4 add_5956_8_lut (.I0(GND_net), .I1(n3369[28]), .I2(n2810), 
            .I3(n17372), .O(n3368[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_8 (.CI(n17372), .I0(n3369[28]), .I1(n2810), .CO(n17373));
    SB_LUT4 add_5956_7_lut (.I0(GND_net), .I1(n3369[27]), .I2(n2810), 
            .I3(n17371), .O(n3368[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_7 (.CI(n17371), .I0(n3369[27]), .I1(n2810), .CO(n17372));
    SB_LUT4 add_5956_6_lut (.I0(GND_net), .I1(n3369[26]), .I2(n2810), 
            .I3(n17370), .O(n3368[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_6 (.CI(n17370), .I0(n3369[26]), .I1(n2810), .CO(n17371));
    SB_LUT4 add_5956_5_lut (.I0(GND_net), .I1(n3369[25]), .I2(n2810), 
            .I3(n17369), .O(n3368[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_5 (.CI(n17369), .I0(n3369[25]), .I1(n2810), .CO(n17370));
    SB_LUT4 add_5956_4_lut (.I0(GND_net), .I1(n3369[24]), .I2(n2810), 
            .I3(n17368), .O(n3368[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_4 (.CI(n17368), .I0(n3369[24]), .I1(n2810), .CO(n17369));
    SB_LUT4 add_5956_3_lut (.I0(GND_net), .I1(n3369[23]), .I2(n2810), 
            .I3(n17367), .O(n3368[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_3 (.CI(n17367), .I0(n3369[23]), .I1(n2810), .CO(n17368));
    SB_LUT4 add_5956_2_lut (.I0(GND_net), .I1(n2813), .I2(GND_net), .I3(GND_net), 
            .O(n3368[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5956_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5956_2 (.CI(GND_net), .I0(n2813), .I1(GND_net), .CO(n17367));
    SB_LUT4 add_5955_10_lut (.I0(GND_net), .I1(n3368[30]), .I2(GND_net), 
            .I3(n17365), .O(n3367[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5955_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5955_10 (.CI(n17365), .I0(n3368[30]), .I1(GND_net), .CO(n3212));
    SB_LUT4 add_5955_9_lut (.I0(GND_net), .I1(n3368[29]), .I2(n2807), 
            .I3(n17364), .O(n3367[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5955_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5955_9 (.CI(n17364), .I0(n3368[29]), .I1(n2807), .CO(n17365));
    SB_LUT4 add_5955_8_lut (.I0(GND_net), .I1(n3368[28]), .I2(n2807), 
            .I3(n17363), .O(n3367[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5955_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5955_8 (.CI(n17363), .I0(n3368[28]), .I1(n2807), .CO(n17364));
    SB_CARRY add_5955_7 (.CI(n17362), .I0(n3368[27]), .I1(n2807), .CO(n17363));
    SB_CARRY add_5955_6 (.CI(n17361), .I0(n3368[26]), .I1(n2807), .CO(n17362));
    SB_CARRY add_5955_5 (.CI(n17360), .I0(n3368[25]), .I1(n2807), .CO(n17361));
    SB_CARRY add_5955_4 (.CI(n17359), .I0(n3368[24]), .I1(n2807), .CO(n17360));
    SB_CARRY add_5955_3 (.CI(n17358), .I0(n3368[23]), .I1(n2807), .CO(n17359));
    SB_CARRY add_5955_2 (.CI(GND_net), .I0(n2810), .I1(GND_net), .CO(n17358));
    SB_LUT4 add_5928_10_lut (.I0(GND_net), .I1(n7546[7]), .I2(n2652), 
            .I3(n17357), .O(n7464[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5928_9_lut (.I0(GND_net), .I1(n7546[6]), .I2(n2652), .I3(n17356), 
            .O(n7464[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_9 (.CI(n17356), .I0(n7546[6]), .I1(n2652), .CO(n17357));
    SB_LUT4 add_5928_8_lut (.I0(GND_net), .I1(n7546[5]), .I2(n2652), .I3(n17355), 
            .O(n7464[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_8 (.CI(n17355), .I0(n7546[5]), .I1(n2652), .CO(n17356));
    SB_LUT4 add_5928_7_lut (.I0(GND_net), .I1(n7546[4]), .I2(n2652), .I3(n17354), 
            .O(n7464[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_7 (.CI(n17354), .I0(n7546[4]), .I1(n2652), .CO(n17355));
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_7 (.CI(n15464), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15465));
    SB_LUT4 add_5928_6_lut (.I0(GND_net), .I1(n7546[3]), .I2(n2652), .I3(n17353), 
            .O(n7464[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_6 (.CI(n17353), .I0(n7546[3]), .I1(n2652), .CO(n17354));
    SB_LUT4 add_5928_5_lut (.I0(GND_net), .I1(n7546[2]), .I2(n2652), .I3(n17352), 
            .O(n7464[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_5 (.CI(n17352), .I0(n7546[2]), .I1(n2652), .CO(n17353));
    SB_LUT4 add_5928_4_lut (.I0(GND_net), .I1(n7546[1]), .I2(n2652), .I3(n17351), 
            .O(n7464[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_4 (.CI(n17351), .I0(n7546[1]), .I1(n2652), .CO(n17352));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15463), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_5928_3_lut (.I0(GND_net), .I1(n7546[0]), .I2(GND_net), 
            .I3(n17350), .O(n7464[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_3 (.CI(n17350), .I0(n7546[0]), .I1(GND_net), .CO(n17351));
    SB_LUT4 add_5928_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2652), .I3(GND_net), .O(n7464[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5928_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5928_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2652), .CO(n17350));
    SB_LUT4 add_6236_8_lut (.I0(GND_net), .I1(n8171[5]), .I2(n2652), .I3(n17349), 
            .O(n7890[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6236_7_lut (.I0(GND_net), .I1(n8171[4]), .I2(n2652), .I3(n17348), 
            .O(n7890[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2831), .I3(GND_net), .O(n3375[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_3 (.CI(n17431), .I0(n3376[22]), 
            .I1(GND_net), .CO(n17432));
    SB_CARRY add_6236_7 (.CI(n17348), .I0(n8171[4]), .I1(n2652), .CO(n17349));
    SB_LUT4 add_6236_6_lut (.I0(GND_net), .I1(n8171[3]), .I2(n2652), .I3(n17347), 
            .O(n7890[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_3_lut (.I0(GND_net), .I1(n3376[22]), 
            .I2(GND_net), .I3(n17431), .O(n3375[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6236_6 (.CI(n17347), .I0(n8171[3]), .I1(n2652), .CO(n17348));
    SB_LUT4 add_6236_5_lut (.I0(GND_net), .I1(n8171[2]), .I2(n2652), .I3(n17346), 
            .O(n7890[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6236_5 (.CI(n17346), .I0(n8171[2]), .I1(n2652), .CO(n17347));
    SB_LUT4 add_6236_4_lut (.I0(GND_net), .I1(n8171[1]), .I2(n2652), .I3(n17345), 
            .O(n7890[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6236_4 (.CI(n17345), .I0(n8171[1]), .I1(n2652), .CO(n17346));
    SB_LUT4 add_6236_3_lut (.I0(GND_net), .I1(n8171[0]), .I2(GND_net), 
            .I3(n17344), .O(n7890[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6236_3 (.CI(n17344), .I0(n8171[0]), .I1(GND_net), .CO(n17345));
    SB_LUT4 add_6236_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2652), .I3(GND_net), .O(n7890[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6236_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6236_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2652), .CO(n17344));
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2831), .CO(n17431));
    SB_LUT4 add_5953_9_lut (.I0(GND_net), .I1(n7890[6]), .I2(n2652), .I3(n17343), 
            .O(n7546[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5953_8_lut (.I0(GND_net), .I1(n7890[5]), .I2(n2652), .I3(n17342), 
            .O(n7546[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_8 (.CI(n17342), .I0(n7890[5]), .I1(n2652), .CO(n17343));
    SB_LUT4 add_5953_7_lut (.I0(GND_net), .I1(n7890[4]), .I2(n2652), .I3(n17341), 
            .O(n7546[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_7 (.CI(n17341), .I0(n7890[4]), .I1(n2652), .CO(n17342));
    SB_LUT4 add_5953_6_lut (.I0(GND_net), .I1(n7890[3]), .I2(n2652), .I3(n17340), 
            .O(n7546[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_6 (.CI(n17340), .I0(n7890[3]), .I1(n2652), .CO(n17341));
    SB_LUT4 add_5953_5_lut (.I0(GND_net), .I1(n7890[2]), .I2(n2652), .I3(n17339), 
            .O(n7546[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_5 (.CI(n17339), .I0(n7890[2]), .I1(n2652), .CO(n17340));
    SB_LUT4 add_5953_4_lut (.I0(GND_net), .I1(n7890[1]), .I2(n2652), .I3(n17338), 
            .O(n7546[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_4 (.CI(n17338), .I0(n7890[1]), .I1(n2652), .CO(n17339));
    SB_LUT4 add_5953_3_lut (.I0(GND_net), .I1(n7890[0]), .I2(GND_net), 
            .I3(n17337), .O(n7546[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_3 (.CI(n17337), .I0(n7890[0]), .I1(GND_net), .CO(n17338));
    SB_LUT4 add_5953_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2652), .I3(GND_net), .O(n7546[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5953_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5953_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2652), .CO(n17337));
    SB_LUT4 add_6484_7_lut (.I0(GND_net), .I1(n8488[3]), .I2(n2652), .I3(n17336), 
            .O(n8171[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6484_6_lut (.I0(GND_net), .I1(n8488[3]), .I2(n2652), .I3(n17335), 
            .O(n8171[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_6 (.CI(n17335), .I0(n8488[3]), .I1(n2652), .CO(n17336));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_4_lut (.I0(GND_net), .I1(n3376[23]), 
            .I2(n2831), .I3(n17432), .O(n3375[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6484_5_lut (.I0(GND_net), .I1(n8488[3]), .I2(n2652), .I3(n17334), 
            .O(n8171[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_5 (.CI(n17334), .I0(n8488[3]), .I1(n2652), .CO(n17335));
    SB_LUT4 add_6484_4_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2652), .I3(n17333), .O(n8171[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_4 (.CI(n17333), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2652), .CO(n17334));
    SB_LUT4 add_6484_3_lut (.I0(GND_net), .I1(n8488[3]), .I2(GND_net), 
            .I3(n17332), .O(n8171[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_3 (.CI(n17332), .I0(n8488[3]), .I1(GND_net), .CO(n17333));
    SB_LUT4 add_6484_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2652), .I3(GND_net), .O(n8171[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6484_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6484_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2652), .CO(n17332));
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_11 (.CI(n17429), .I0(n3375[30]), 
            .I1(GND_net), .CO(n3240));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_10_lut (.I0(GND_net), .I1(n3375[29]), 
            .I2(n2828), .I3(n17428), .O(n3374[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_6 (.CI(n15463), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15464));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(\Amp25_out1[14] ), .I3(n15462), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Look_Up_Table_f1_31__I_0_i1719_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Look_Up_Table_sub_temp1[15]), .I2(GND_net), .I3(GND_net), 
            .O(n2652));   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(378[31:76])
    defparam Look_Up_Table_f1_31__I_0_i1719_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_5 (.CI(n15462), .I0(GND_net), 
            .I1(\Amp25_out1[14] ), .CO(n15463));
    SB_LUT4 Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut (.I0(\Product_mul_temp[26] ), 
            .I1(GND_net), .I2(VCC_net), .I3(n15461), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_sub_temp1_15__I_0_add_2_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3098_17_lut (.I0(GND_net), .I1(n3380[31]), .I2(n3260), 
            .I3(n17504), .O(Look_Up_Table_mul_temp1[47])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_16_lut (.I0(GND_net), .I1(n3379[31]), .I2(n3256), 
            .I3(n17503), .O(Look_Up_Table_mul_temp1[46])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_16 (.CI(n17503), .I0(n3379[31]), .I1(n3256), .CO(n17504));
    SB_LUT4 add_3098_15_lut (.I0(GND_net), .I1(n3378[31]), .I2(n3252), 
            .I3(n17502), .O(Look_Up_Table_mul_temp1[45])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_15 (.CI(n17502), .I0(n3378[31]), .I1(n3252), .CO(n17503));
    SB_LUT4 add_3098_14_lut (.I0(GND_net), .I1(n3377[31]), .I2(n3248), 
            .I3(n17501), .O(Look_Up_Table_mul_temp1[44])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_14 (.CI(n17501), .I0(n3377[31]), .I1(n3248), .CO(n17502));
    SB_LUT4 add_3098_13_lut (.I0(GND_net), .I1(n3376[31]), .I2(n3244), 
            .I3(n17500), .O(Look_Up_Table_mul_temp1[43])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_13 (.CI(n17500), .I0(n3376[31]), .I1(n3244), .CO(n17501));
    SB_LUT4 add_3098_12_lut (.I0(GND_net), .I1(n3375[31]), .I2(n3240), 
            .I3(n17499), .O(Look_Up_Table_mul_temp1[42])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_12 (.CI(n17499), .I0(n3375[31]), .I1(n3240), .CO(n17500));
    SB_LUT4 add_3098_11_lut (.I0(GND_net), .I1(n3374[31]), .I2(n3236), 
            .I3(n17498), .O(Look_Up_Table_mul_temp1[41])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_11 (.CI(n17498), .I0(n3374[31]), .I1(n3236), .CO(n17499));
    SB_LUT4 add_3098_10_lut (.I0(GND_net), .I1(n3373[31]), .I2(n3232), 
            .I3(n17497), .O(Look_Up_Table_mul_temp1[40])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_10 (.CI(n17497), .I0(n3373[31]), .I1(n3232), .CO(n17498));
    SB_LUT4 add_3098_9_lut (.I0(GND_net), .I1(n3372[31]), .I2(n3228), 
            .I3(n17496), .O(Look_Up_Table_mul_temp1[39])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_9 (.CI(n17496), .I0(n3372[31]), .I1(n3228), .CO(n17497));
    SB_LUT4 add_3098_8_lut (.I0(GND_net), .I1(n3371[31]), .I2(n3224), 
            .I3(n17495), .O(Look_Up_Table_mul_temp1[38])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_8 (.CI(n17495), .I0(n3371[31]), .I1(n3224), .CO(n17496));
    SB_LUT4 add_3098_7_lut (.I0(GND_net), .I1(n3370[31]), .I2(n3220), 
            .I3(n17494), .O(Look_Up_Table_mul_temp1[37])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_7 (.CI(n17494), .I0(n3370[31]), .I1(n3220), .CO(n17495));
    SB_LUT4 add_3098_6_lut (.I0(GND_net), .I1(n3369[31]), .I2(n3216), 
            .I3(n17493), .O(Look_Up_Table_mul_temp1[36])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_6 (.CI(n17493), .I0(n3369[31]), .I1(n3216), .CO(n17494));
    SB_LUT4 add_3098_5_lut (.I0(GND_net), .I1(n3368[31]), .I2(n3212), 
            .I3(n17492), .O(Look_Up_Table_mul_temp1[35])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_5 (.CI(n17492), .I0(n3368[31]), .I1(n3212), .CO(n17493));
    SB_LUT4 add_3098_4_lut (.I0(GND_net), .I1(n3367[31]), .I2(GND_net), 
            .I3(n17491), .O(Look_Up_Table_mul_temp1[34])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_4 (.CI(n17491), .I0(n3367[31]), .I1(GND_net), .CO(n17492));
    SB_LUT4 add_3098_3_lut (.I0(GND_net), .I1(n3367[30]), .I2(GND_net), 
            .I3(n17490), .O(Look_Up_Table_out1_1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_3 (.CI(n17490), .I0(n3367[30]), .I1(GND_net), .CO(n17491));
    SB_LUT4 add_3098_2_lut (.I0(GND_net), .I1(n3367[29]), .I2(Look_Up_Table_sub_temp1[15]), 
            .I3(GND_net), .O(Look_Up_Table_out1_1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_2 (.CI(GND_net), .I0(n3367[29]), .I1(Look_Up_Table_sub_temp1[15]), 
            .CO(n17490));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_11_lut (.I0(GND_net), .I1(n7464[8]), 
            .I2(GND_net), .I3(n17489), .O(n3380[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_10_lut (.I0(GND_net), .I1(n7464[7]), 
            .I2(n2652), .I3(n17488), .O(n3380[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_10 (.CI(n17488), .I0(n7464[7]), 
            .I1(n2652), .CO(n17489));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_9_lut (.I0(GND_net), .I1(n7464[6]), 
            .I2(n2652), .I3(n17487), .O(n3380[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_9 (.CI(n17487), .I0(n7464[6]), 
            .I1(n2652), .CO(n17488));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_8_lut (.I0(GND_net), .I1(n7464[5]), 
            .I2(n2652), .I3(n17486), .O(n3380[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_8 (.CI(n17486), .I0(n7464[5]), 
            .I1(n2652), .CO(n17487));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_7_lut (.I0(GND_net), .I1(n7464[4]), 
            .I2(n2652), .I3(n17485), .O(n3380[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_7 (.CI(n17485), .I0(n7464[4]), 
            .I1(n2652), .CO(n17486));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_6_lut (.I0(GND_net), .I1(n7464[3]), 
            .I2(n2652), .I3(n17484), .O(n3380[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_6 (.CI(n17484), .I0(n7464[3]), 
            .I1(n2652), .CO(n17485));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_5_lut (.I0(GND_net), .I1(n7464[2]), 
            .I2(n2652), .I3(n17483), .O(n3380[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_5 (.CI(n17483), .I0(n7464[2]), 
            .I1(n2652), .CO(n17484));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_4_lut (.I0(GND_net), .I1(n7464[1]), 
            .I2(n2652), .I3(n17482), .O(n3380[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_4 (.CI(n17482), .I0(n7464[1]), 
            .I1(n2652), .CO(n17483));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_3_lut (.I0(GND_net), .I1(n7464[0]), 
            .I2(GND_net), .I3(n17481), .O(n3380[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_3 (.CI(n17481), .I0(n7464[0]), 
            .I1(GND_net), .CO(n17482));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2276_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2652), .I3(GND_net), .O(n3380[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2276_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2276_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2652), .CO(n17481));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_11_lut (.I0(GND_net), .I1(n3380[30]), 
            .I2(GND_net), .I3(n17479), .O(n3379[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_11 (.CI(n17479), .I0(n3380[30]), 
            .I1(GND_net), .CO(n3260));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_10_lut (.I0(GND_net), .I1(n3380[29]), 
            .I2(n2843), .I3(n17478), .O(n3379[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_10 (.CI(n17478), .I0(n3380[29]), 
            .I1(n2843), .CO(n17479));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_9_lut (.I0(GND_net), .I1(n3380[28]), 
            .I2(n2843), .I3(n17477), .O(n3379[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_9 (.CI(n17477), .I0(n3380[28]), 
            .I1(n2843), .CO(n17478));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_8_lut (.I0(GND_net), .I1(n3380[27]), 
            .I2(n2843), .I3(n17476), .O(n3379[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_8 (.CI(n17476), .I0(n3380[27]), 
            .I1(n2843), .CO(n17477));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_7_lut (.I0(GND_net), .I1(n3380[26]), 
            .I2(n2843), .I3(n17475), .O(n3379[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_7 (.CI(n17475), .I0(n3380[26]), 
            .I1(n2843), .CO(n17476));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_6_lut (.I0(GND_net), .I1(n3380[25]), 
            .I2(n2843), .I3(n17474), .O(n3379[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_6 (.CI(n17474), .I0(n3380[25]), 
            .I1(n2843), .CO(n17475));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_5_lut (.I0(GND_net), .I1(n3380[24]), 
            .I2(n2843), .I3(n17473), .O(n3379[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_5 (.CI(n17473), .I0(n3380[24]), 
            .I1(n2843), .CO(n17474));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_4_lut (.I0(GND_net), .I1(n3380[23]), 
            .I2(n2843), .I3(n17472), .O(n3379[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_4 (.CI(n17472), .I0(n3380[23]), 
            .I1(n2843), .CO(n17473));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_3_lut (.I0(GND_net), .I1(n3380[22]), 
            .I2(GND_net), .I3(n17471), .O(n3379[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_3 (.CI(n17471), .I0(n3380[22]), 
            .I1(GND_net), .CO(n17472));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2275_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2843), .I3(GND_net), .O(n3379[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2275_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2275_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2843), .CO(n17471));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_11_lut (.I0(GND_net), .I1(n3379[30]), 
            .I2(GND_net), .I3(n17469), .O(n3378[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_11 (.CI(n17469), .I0(n3379[30]), 
            .I1(GND_net), .CO(n3256));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_10_lut (.I0(GND_net), .I1(n3379[29]), 
            .I2(n2840), .I3(n17468), .O(n3378[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_10 (.CI(n17468), .I0(n3379[29]), 
            .I1(n2840), .CO(n17469));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_9_lut (.I0(GND_net), .I1(n3379[28]), 
            .I2(n2840), .I3(n17467), .O(n3378[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_9 (.CI(n17467), .I0(n3379[28]), 
            .I1(n2840), .CO(n17468));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_8_lut (.I0(GND_net), .I1(n3379[27]), 
            .I2(n2840), .I3(n17466), .O(n3378[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_8 (.CI(n17466), .I0(n3379[27]), 
            .I1(n2840), .CO(n17467));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_7_lut (.I0(GND_net), .I1(n3379[26]), 
            .I2(n2840), .I3(n17465), .O(n3378[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_7 (.CI(n17465), .I0(n3379[26]), 
            .I1(n2840), .CO(n17466));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_6_lut (.I0(GND_net), .I1(n3379[25]), 
            .I2(n2840), .I3(n17464), .O(n3378[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_6 (.CI(n17464), .I0(n3379[25]), 
            .I1(n2840), .CO(n17465));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_5_lut (.I0(GND_net), .I1(n3379[24]), 
            .I2(n2840), .I3(n17463), .O(n3378[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_5 (.CI(n17463), .I0(n3379[24]), 
            .I1(n2840), .CO(n17464));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_4_lut (.I0(GND_net), .I1(n3379[23]), 
            .I2(n2840), .I3(n17462), .O(n3378[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_4 (.CI(n17462), .I0(n3379[23]), 
            .I1(n2840), .CO(n17463));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_3_lut (.I0(GND_net), .I1(n3379[22]), 
            .I2(GND_net), .I3(n17461), .O(n3378[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_3 (.CI(n17461), .I0(n3379[22]), 
            .I1(GND_net), .CO(n17462));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2274_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2840), .I3(GND_net), .O(n3378[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2274_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2274_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2840), .CO(n17461));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_11_lut (.I0(GND_net), .I1(n3378[30]), 
            .I2(GND_net), .I3(n17459), .O(n3377[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_11 (.CI(n17459), .I0(n3378[30]), 
            .I1(GND_net), .CO(n3252));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_10_lut (.I0(GND_net), .I1(n3378[29]), 
            .I2(n2840), .I3(n17458), .O(n3377[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_10 (.CI(n17458), .I0(n3378[29]), 
            .I1(n2840), .CO(n17459));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_9_lut (.I0(GND_net), .I1(n3378[28]), 
            .I2(n2840), .I3(n17457), .O(n3377[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_9 (.CI(n17457), .I0(n3378[28]), 
            .I1(n2840), .CO(n17458));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_8_lut (.I0(GND_net), .I1(n3378[27]), 
            .I2(n2840), .I3(n17456), .O(n3377[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_8 (.CI(n17456), .I0(n3378[27]), 
            .I1(n2840), .CO(n17457));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_7_lut (.I0(GND_net), .I1(n3378[26]), 
            .I2(n2840), .I3(n17455), .O(n3377[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_7 (.CI(n17455), .I0(n3378[26]), 
            .I1(n2840), .CO(n17456));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_6_lut (.I0(GND_net), .I1(n3378[25]), 
            .I2(n2840), .I3(n17454), .O(n3377[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_6 (.CI(n17454), .I0(n3378[25]), 
            .I1(n2840), .CO(n17455));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_5_lut (.I0(GND_net), .I1(n3378[24]), 
            .I2(n2840), .I3(n17453), .O(n3377[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_5 (.CI(n17453), .I0(n3378[24]), 
            .I1(n2840), .CO(n17454));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_4_lut (.I0(GND_net), .I1(n3378[23]), 
            .I2(n2840), .I3(n17452), .O(n3377[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_4 (.CI(n17452), .I0(n3378[23]), 
            .I1(n2840), .CO(n17453));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_3_lut (.I0(GND_net), .I1(n3378[22]), 
            .I2(GND_net), .I3(n17451), .O(n3377[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_3 (.CI(n17451), .I0(n3378[22]), 
            .I1(GND_net), .CO(n17452));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2273_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2840), .I3(GND_net), .O(n3377[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2273_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2273_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2840), .CO(n17451));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_11_lut (.I0(GND_net), .I1(n3377[30]), 
            .I2(GND_net), .I3(n17449), .O(n3376[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_11 (.CI(n17449), .I0(n3377[30]), 
            .I1(GND_net), .CO(n3248));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_10_lut (.I0(GND_net), .I1(n3377[29]), 
            .I2(n2834), .I3(n17448), .O(n3376[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_10 (.CI(n17448), .I0(n3377[29]), 
            .I1(n2834), .CO(n17449));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_9_lut (.I0(GND_net), .I1(n3377[28]), 
            .I2(n2834), .I3(n17447), .O(n3376[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_9 (.CI(n17447), .I0(n3377[28]), 
            .I1(n2834), .CO(n17448));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_8_lut (.I0(GND_net), .I1(n3377[27]), 
            .I2(n2834), .I3(n17446), .O(n3376[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_8 (.CI(n17446), .I0(n3377[27]), 
            .I1(n2834), .CO(n17447));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_7_lut (.I0(GND_net), .I1(n3377[26]), 
            .I2(n2834), .I3(n17445), .O(n3376[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_7 (.CI(n17445), .I0(n3377[26]), 
            .I1(n2834), .CO(n17446));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_6_lut (.I0(GND_net), .I1(n3377[25]), 
            .I2(n2834), .I3(n17444), .O(n3376[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_6 (.CI(n17444), .I0(n3377[25]), 
            .I1(n2834), .CO(n17445));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_5_lut (.I0(GND_net), .I1(n3377[24]), 
            .I2(n2834), .I3(n17443), .O(n3376[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_5 (.CI(n17443), .I0(n3377[24]), 
            .I1(n2834), .CO(n17444));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_4_lut (.I0(GND_net), .I1(n3377[23]), 
            .I2(n2834), .I3(n17442), .O(n3376[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_4 (.CI(n17442), .I0(n3377[23]), 
            .I1(n2834), .CO(n17443));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_3_lut (.I0(GND_net), .I1(n3377[22]), 
            .I2(GND_net), .I3(n17441), .O(n3376[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_3 (.CI(n17441), .I0(n3377[22]), 
            .I1(GND_net), .CO(n17442));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2272_2_lut (.I0(GND_net), .I1(Look_Up_Table_sub_temp1[15]), 
            .I2(n2834), .I3(GND_net), .O(n3376[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2272_2 (.CI(GND_net), .I0(Look_Up_Table_sub_temp1[15]), 
            .I1(n2834), .CO(n17441));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_11_lut (.I0(GND_net), .I1(n3376[30]), 
            .I2(GND_net), .I3(n17439), .O(n3375[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_11 (.CI(n17439), .I0(n3376[30]), 
            .I1(GND_net), .CO(n3244));
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_10 (.CI(n17428), .I0(n3375[29]), 
            .I1(n2828), .CO(n17429));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_9_lut (.I0(GND_net), .I1(n3375[28]), 
            .I2(n2828), .I3(n17427), .O(n3374[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_9 (.CI(n17427), .I0(n3375[28]), 
            .I1(n2828), .CO(n17428));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_8_lut (.I0(GND_net), .I1(n3375[27]), 
            .I2(n2828), .I3(n17426), .O(n3374[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_8 (.CI(n17426), .I0(n3375[27]), 
            .I1(n2828), .CO(n17427));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_7_lut (.I0(GND_net), .I1(n3375[26]), 
            .I2(n2828), .I3(n17425), .O(n3374[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_10_lut (.I0(GND_net), .I1(n3376[29]), 
            .I2(n2831), .I3(n17438), .O(n3375[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_7 (.CI(n17425), .I0(n3375[26]), 
            .I1(n2828), .CO(n17426));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_6_lut (.I0(GND_net), .I1(n3375[25]), 
            .I2(n2828), .I3(n17424), .O(n3374[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_10 (.CI(n17438), .I0(n3376[29]), 
            .I1(n2831), .CO(n17439));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_9_lut (.I0(GND_net), .I1(n3376[28]), 
            .I2(n2831), .I3(n17437), .O(n3375[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_sub_temp1_15__I_0_add_2_4 (.CI(n15461), .I0(GND_net), 
            .I1(VCC_net), .CO(n15462));
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2270_6 (.CI(n17424), .I0(n3375[25]), 
            .I1(n2828), .CO(n17425));
    SB_LUT4 add_551_15_lut (.I0(GND_net), .I1(GND_net), .I2(Look_Up_Table_mul_temp1[47]), 
            .I3(n15956), .O(Look_Up_Table_out1_1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_551_14_lut (.I0(GND_net), .I1(\Amp25_out1[14] ), .I2(Look_Up_Table_mul_temp1[46]), 
            .I3(n15955), .O(Look_Up_Table_out1_1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_14 (.CI(n15955), .I0(\Amp25_out1[14] ), .I1(Look_Up_Table_mul_temp1[46]), 
            .CO(n15956));
    SB_LUT4 add_551_13_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[45]), 
            .I3(n15954), .O(Look_Up_Table_out1_1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_13 (.CI(n15954), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[45]), 
            .CO(n15955));
    SB_LUT4 add_551_12_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[44]), 
            .I3(n15953), .O(Look_Up_Table_out1_1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_12 (.CI(n15953), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[44]), 
            .CO(n15954));
    SB_LUT4 add_551_11_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[43]), 
            .I3(n15952), .O(Look_Up_Table_out1_1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_11 (.CI(n15952), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[43]), 
            .CO(n15953));
    SB_LUT4 add_551_10_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[42]), 
            .I3(n15951), .O(Look_Up_Table_out1_1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_10 (.CI(n15951), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[42]), 
            .CO(n15952));
    SB_LUT4 add_551_9_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[41]), 
            .I3(n15950), .O(Look_Up_Table_out1_1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_9 (.CI(n15950), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[41]), 
            .CO(n15951));
    SB_LUT4 add_551_8_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[40]), 
            .I3(n15949), .O(Look_Up_Table_out1_1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_8 (.CI(n15949), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[40]), 
            .CO(n15950));
    SB_LUT4 add_551_7_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[39]), 
            .I3(n15948), .O(Look_Up_Table_out1_1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_7 (.CI(n15948), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[39]), 
            .CO(n15949));
    SB_LUT4 add_551_6_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[38]), 
            .I3(n15947), .O(Look_Up_Table_out1_1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_6 (.CI(n15947), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[38]), 
            .CO(n15948));
    SB_LUT4 add_551_5_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[37]), 
            .I3(n15946), .O(Look_Up_Table_out1_1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_5 (.CI(n15946), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[37]), 
            .CO(n15947));
    SB_LUT4 add_551_4_lut (.I0(GND_net), .I1(GND_net), .I2(Look_Up_Table_mul_temp1[36]), 
            .I3(n15945), .O(Look_Up_Table_out1_1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_4 (.CI(n15945), .I0(GND_net), .I1(Look_Up_Table_mul_temp1[36]), 
            .CO(n15946));
    SB_LUT4 add_551_3_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[35]), 
            .I3(n15944), .O(Look_Up_Table_out1_1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_3 (.CI(n15944), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[35]), 
            .CO(n15945));
    SB_LUT4 add_551_2_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_mul_temp1[34]), 
            .I3(GND_net), .O(Look_Up_Table_out1_1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_551_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_551_2 (.CI(GND_net), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_mul_temp1[34]), 
            .CO(n15944));
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_9 (.CI(n17437), .I0(n3376[28]), 
            .I1(n2831), .CO(n17438));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_8_lut (.I0(GND_net), .I1(n3376[27]), 
            .I2(n2831), .I3(n17436), .O(n3375[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_8 (.CI(n17436), .I0(n3376[27]), 
            .I1(n2831), .CO(n17437));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2270_5_lut (.I0(GND_net), .I1(n3375[24]), 
            .I2(n2828), .I3(n17423), .O(n3374[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2270_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_7_lut (.I0(GND_net), .I1(n3376[26]), 
            .I2(n2831), .I3(n17435), .O(n3375[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_7 (.CI(n17435), .I0(n3376[26]), 
            .I1(n2831), .CO(n17436));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_6_lut (.I0(GND_net), .I1(n3376[25]), 
            .I2(n2831), .I3(n17434), .O(n3375[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_6 (.CI(n17434), .I0(n3376[25]), 
            .I1(n2831), .CO(n17435));
    SB_LUT4 Look_Up_Table_f1_31__I_0_add_2271_5_lut (.I0(GND_net), .I1(n3376[24]), 
            .I2(n2831), .I3(n17433), .O(n3375[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Look_Up_Table_f1_31__I_0_add_2271_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Look_Up_Table_f1_31__I_0_add_2271_5 (.CI(n17433), .I0(n3376[24]), 
            .I1(n2831), .CO(n17434));
    SB_LUT4 u_29__I_0_71_inv_0_i4_1_lut (.I0(\Product_mul_temp[26] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\Amp25_out1[14] ));   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(281[23:56])
    defparam u_29__I_0_71_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13555_2_lut (.I0(Look_Up_Table_sub_temp1[15]), .I1(\Amp25_out1[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n8488[3]));   // ../../hdlcoderFocCurrentFixptHdl/Sine_Cosine_LUT.v(378[31:76])
    defparam i13555_2_lut.LUT_INIT = 16'h8888;
    VCC i1 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module Park_Transform
//

module Park_Transform (GND_net, n628, n142, \Product_mul_temp[26] , 
            Look_Up_Table_out1_1, \dCurrent[31] , \dCurrent[30] , \dCurrent[29] , 
            \dCurrent[28] , \dCurrent[27] , \dCurrent[26] , \dCurrent[25] , 
            \dCurrent[24] , \dCurrent[23] , \dCurrent[22] , \dCurrent[21] , 
            \dCurrent[20] , \dCurrent[19] , \dCurrent[18] , \dCurrent[17] , 
            \dCurrent[16] , \dCurrent[15] , \dCurrent[14] , \dCurrent[13] , 
            \dCurrent[12] , \dCurrent[11] , \dCurrent[10] , \dCurrent[9] , 
            \dCurrent[8] , \dCurrent[7] , \dCurrent[6] , \dCurrent[5] , 
            \dCurrent[4] , \qCurrent[3] , \dCurrent[3] , n139, n794, 
            \qCurrent[31] , \qCurrent[30] , \qCurrent[29] , \qCurrent[28] , 
            \qCurrent[27] , \qCurrent[26] , \qCurrent[25] , \qCurrent[24] , 
            \qCurrent[23] , \qCurrent[22] , \qCurrent[21] , \qCurrent[20] , 
            \qCurrent[19] , \qCurrent[18] , \qCurrent[17] , \qCurrent[16] , 
            \qCurrent[15] , \qCurrent[14] , \qCurrent[13] , \qCurrent[12] , 
            \qCurrent[11] , \qCurrent[10] , \qCurrent[9] , \qCurrent[8] , 
            \qCurrent[7] , \qCurrent[6] , \qCurrent[5] , \qCurrent[4] , 
            \Amp25_out1[14] , n4) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n628;
    input n142;
    input \Product_mul_temp[26] ;
    input [15:0]Look_Up_Table_out1_1;
    output \dCurrent[31] ;
    output \dCurrent[30] ;
    output \dCurrent[29] ;
    output \dCurrent[28] ;
    output \dCurrent[27] ;
    output \dCurrent[26] ;
    output \dCurrent[25] ;
    output \dCurrent[24] ;
    output \dCurrent[23] ;
    output \dCurrent[22] ;
    output \dCurrent[21] ;
    output \dCurrent[20] ;
    output \dCurrent[19] ;
    output \dCurrent[18] ;
    output \dCurrent[17] ;
    output \dCurrent[16] ;
    output \dCurrent[15] ;
    output \dCurrent[14] ;
    output \dCurrent[13] ;
    output \dCurrent[12] ;
    output \dCurrent[11] ;
    output \dCurrent[10] ;
    output \dCurrent[9] ;
    output \dCurrent[8] ;
    output \dCurrent[7] ;
    output \dCurrent[6] ;
    output \dCurrent[5] ;
    output \dCurrent[4] ;
    output \qCurrent[3] ;
    output \dCurrent[3] ;
    input n139;
    input n794;
    output \qCurrent[31] ;
    output \qCurrent[30] ;
    output \qCurrent[29] ;
    output \qCurrent[28] ;
    output \qCurrent[27] ;
    output \qCurrent[26] ;
    output \qCurrent[25] ;
    output \qCurrent[24] ;
    output \qCurrent[23] ;
    output \qCurrent[22] ;
    output \qCurrent[21] ;
    output \qCurrent[20] ;
    output \qCurrent[19] ;
    output \qCurrent[18] ;
    output \qCurrent[17] ;
    output \qCurrent[16] ;
    output \qCurrent[15] ;
    output \qCurrent[14] ;
    output \qCurrent[13] ;
    output \qCurrent[12] ;
    output \qCurrent[11] ;
    output \qCurrent[10] ;
    output \qCurrent[9] ;
    output \qCurrent[8] ;
    output \qCurrent[7] ;
    output \qCurrent[6] ;
    output \qCurrent[5] ;
    output \qCurrent[4] ;
    input \Amp25_out1[14] ;
    input n4;
    
    
    wire n17184;
    wire [14:0]n838;
    
    wire n604, n17185;
    wire [14:0]n837;
    
    wire n17183;
    wire [14:0]n840;
    wire [14:0]n841;
    
    wire n769, n16961, n17034;
    wire [14:0]n836;
    
    wire n598, n17035, n12, n14, n4_c, n18, n19845, n771;
    wire [14:0]n833;
    wire [14:0]n834;
    
    wire n592, n17058;
    wire [14:0]n839;
    
    wire n610, n16972;
    wire [14:0]n838_adj_2170;
    
    wire n607, n16987, n16988, n17182, n17000, n17001;
    wire [31:0]Product1_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(38[22:39])
    wire [14:0]n835;
    
    wire n747, n17086, n26, n7, n791, n17181;
    wire [14:0]n837_adj_2171;
    
    wire n601, n17012, n17180;
    wire [14:0]n835_adj_2172;
    
    wire n17033, n17179, n17059, n17087, n17178, n17057, n17177, 
        n17176;
    wire [14:0]n834_adj_2173;
    
    wire n743, n17085, n17013, n17032;
    wire [14:0]n842;
    
    wire n773, n16946;
    wire [31:0]Product4_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(43[22:39])
    
    wire n16900, n16901;
    wire [14:0]n845;
    
    wire n785;
    wire [14:0]n839_adj_2174;
    
    wire n761, n17174, n763;
    wire [14:0]n833_adj_2175;
    
    wire n739, n17084, n17031, n613, n16960, n17030, n16973, n17173, 
        n16986, n16999, n17029, n17028, n17011, n17027, n17083, 
        n17056, n17172, n17026, n17171, n16932;
    wire [14:0]n843;
    
    wire n619, n16933, n17170;
    wire [14:0]n832;
    
    wire n17055;
    wire [14:0]n832_adj_2176;
    
    wire n737, n17081, n17169, n739_adj_2006, n17054, n779, n16911, 
        n16971, n16985, n17053, n17168, n16998, n17167, n17025;
    wire [31:0]dCurrent;   // ../../hdlcoderFocCurrentFixptHdl/FOC_Current_Control.v(78[22:30])
    
    wire n17080, n595, n17024, n17079, n17166, n16959, n745, n17051, 
        n747_adj_2012;
    wire [14:0]n844;
    
    wire n622, n16921, n17165, n17050, n16931, n17078, n17164, 
        n16922, n17163, n16912, n775, n16910, n16920, n16930, 
        n616, n16945, n17162, n16984, n17010, n17023, n17161, 
        n17049;
    wire [14:0]n840_adj_2177;
    
    wire n765, n17159, n767, n16958, n16929, n17158, n17157, n17156, 
        n16909, n17155, n16944, n17154, n16970, n16957, n16983, 
        n16997, n17153, n17048, n17077, n17152, n16996, n17151, 
        n17150, n17149, n17076, n16919, n16928, n16943, n16956, 
        n17148, n16969, n16982, n17009, n17147, n17047, n17046, 
        n17045, n17146, n17044, n16995;
    wire [14:0]n841_adj_2178;
    
    wire n17144, n771_adj_2032, n17075, n17143, n17043, n17142, 
        n16955, n17008, n17074, n17141, n17073, n16942, n753, 
        n17021, n17140, n17072, n16968, n16994, n17139, n17138, 
        n17137, n16981, n16941, n17136, n17135, n17134, n17133, 
        n767_adj_2041, n16908, n16918, n17132, n16927, n16954, n16967, 
        n17131, n757, n17006, n755, n17042, n17071;
    wire [14:0]n842_adj_2179;
    
    wire n17129, n775_adj_2047, n17070, n17020, n17303, n17302, 
        n17301, n17300, n17299, n17298, n17297, n17128, n17296, 
        n16980, n16940, n17295, n17127, n17041, n16917, n17294, 
        n16966, n17126, n16979, n17293, n17292, n17125, n17291, 
        n17290, n763_adj_2054, n16907, n17124, n17123, n16939, n16926, 
        n16938, n16993, n17289, n759, n16953, n17288, n17122, 
        n16952, n16965, n16978, n17019, n17287, n17121, n17005, 
        n17018, n17286, n17069, n17120, n17285, n17119, n17284, 
        n17283, n17282, n17281, n17280, n17040, n17279, n17278, 
        n16991, n17277, n17004, n17118, n17017, n17039, n17068;
    wire [14:0]n843_adj_2180;
    
    wire n777, n17116, n779_adj_2070, n17264, n17263, n17115, n17262, 
        n17261, n16906, n16916, n16937, n17260, n17114, n17003, 
        n17113, n17259, n17112, n17258, n17257, n17256, n17255, 
        n17254, n17038, n741, n17066, n17111, n16905, n16915, 
        n17253, n16925, n16951, n17110, n16964, n16976, n16990, 
        n17252, n17016, n17109, n17251, n743_adj_2096, n17249, n17248, 
        n17247, n17246, n17065, n17108, n17245, n749, n17244, 
        n17107, n625, n751, n16904, n16936, n17243, n16950, n16975, 
        n781, n16989, n17002, n17015, n17242;
    wire [14:0]n844_adj_2181;
    
    wire n17105, n783, n17241, n17104, n17240, n17239, n17238, 
        n17237, n17064, n17236, n17103, n16903, n16924, n16935, 
        n17234, n17102, n16963, n16974, n17014, n17233, n17101, 
        n17036, n17063, n17100, n17099, n17232, n17231, n17230, 
        n17229, n17228, n17227, n17226, n17225, n17224, n17223, 
        n17098, n17222, n18165, n787, n18164, n18163, n18162, 
        n18161, n18160, n17221;
    wire [14:0]n836_adj_2182;
    
    wire n17219, n751_adj_2142, n16902, n17218, n17217, n17216, 
        n17097, n16949, n17215, n17214, n787_adj_2149, n17096, n17213, 
        n17212, n16914, n17095, n17211, n17210, n17094, n16913, 
        n17209, n17093, n17208, n17092, n17091, n17207, n17206, 
        n17204, n755_adj_2161, n17203, n17202, n17201, n17200, n17199, 
        n17090, n17062, n17198, n759_adj_2166, n17089, n17197, n783_adj_2167, 
        n16948, n17196, n17985, n17984, n17983, n17982, n17981, 
        n17980, n17061, n17195, n17060, n17194, n17193, n17192, 
        n17088, n17191, n17189, n17188, n17187, n17186, VCC_net, 
        n15774, n15773, n15772, n15771, n15770, n15769, n15768, 
        n15767, n15766, n15765, n15764, n15763, n15762, n15761, 
        n15760, n15759, n15758, n15757, n15756, n15755, n15754, 
        n15753, n15752, n15751, n15750, n15749, n15748, n6;
    
    SB_CARRY Alpha_15__I_0_11_add_566_11 (.CI(n17184), .I0(n838[8]), .I1(n604), 
            .CO(n17185));
    SB_LUT4 Alpha_15__I_0_11_add_566_10_lut (.I0(GND_net), .I1(n838[7]), 
            .I2(n604), .I3(n17183), .O(n837[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_16_lut (.I0(GND_net), .I1(n841[11]), .I2(n769), 
            .I3(n16961), .O(n840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_14 (.CI(n17034), .I0(n836[11]), .I1(n598), 
            .CO(n17035));
    SB_LUT4 i1_4_lut (.I0(n628), .I1(n142), .I2(n12), .I3(n14), .O(n4_c));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_4_lut.LUT_INIT = 16'heca8;
    SB_LUT4 i1_4_lut_adj_305 (.I0(n628), .I1(n142), .I2(n14), .I3(n12), 
            .O(n18));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_4_lut_adj_305.LUT_INIT = 16'heca8;
    SB_LUT4 i2_4_lut (.I0(n142), .I1(n4_c), .I2(n628), .I3(n12), .O(n19845));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i2_4_lut.LUT_INIT = 16'heeec;
    SB_CARRY Beta_15__I_0_add_569_16 (.CI(n16961), .I0(n841[11]), .I1(n769), 
            .CO(n771));
    SB_LUT4 Beta_15__I_0_add_562_8_lut (.I0(GND_net), .I1(n834[5]), .I2(n592), 
            .I3(n17058), .O(n833[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_12_lut (.I0(GND_net), .I1(n840[9]), .I2(n610), 
            .I3(n16972), .O(n839[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_12_lut (.I0(GND_net), .I1(n839[9]), .I2(n607), 
            .I3(n16987), .O(n838_adj_2170[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_12 (.CI(n16987), .I0(n839[9]), .I1(n607), 
            .CO(n16988));
    SB_CARRY Alpha_15__I_0_11_add_566_10 (.CI(n17183), .I0(n838[7]), .I1(n604), 
            .CO(n17184));
    SB_LUT4 Alpha_15__I_0_11_add_566_9_lut (.I0(GND_net), .I1(n838[6]), 
            .I2(n604), .I3(n17182), .O(n837[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_9 (.CI(n17182), .I0(n838[6]), .I1(n604), 
            .CO(n17183));
    SB_CARRY Beta_15__I_0_add_566_10 (.CI(n17000), .I0(n838_adj_2170[7]), 
            .I1(n604), .CO(n17001));
    SB_LUT4 add_1234_5_lut (.I0(GND_net), .I1(n835[14]), .I2(n747), .I3(n17086), 
            .O(Product1_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_306 (.I0(n628), .I1(n142), .I2(n19845), .I3(n18), 
            .O(n26));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_4_lut_adj_306.LUT_INIT = 16'heca8;
    SB_LUT4 i1_3_lut (.I0(n142), .I1(n26), .I2(\Product_mul_temp[26] ), 
            .I3(GND_net), .O(n7));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_307 (.I0(n628), .I1(n7), .I2(Look_Up_Table_out1_1[13]), 
            .I3(n26), .O(n791));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_4_lut_adj_307.LUT_INIT = 16'hcecc;
    SB_LUT4 Alpha_15__I_0_11_add_566_8_lut (.I0(GND_net), .I1(n838[5]), 
            .I2(n604), .I3(n17181), .O(n837[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_8 (.CI(n17181), .I0(n838[5]), .I1(n604), 
            .CO(n17182));
    SB_LUT4 Beta_15__I_0_add_565_7_lut (.I0(GND_net), .I1(n837_adj_2171[4]), 
            .I2(n601), .I3(n17012), .O(n836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_566_7_lut (.I0(GND_net), .I1(n838[4]), 
            .I2(n604), .I3(n17180), .O(n837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_13_lut (.I0(GND_net), .I1(n836[10]), .I2(n598), 
            .I3(n17033), .O(n835_adj_2172[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_13 (.CI(n17033), .I0(n836[10]), .I1(n598), 
            .CO(n17034));
    SB_CARRY Alpha_15__I_0_11_add_566_7 (.CI(n17180), .I0(n838[4]), .I1(n604), 
            .CO(n17181));
    SB_LUT4 Alpha_15__I_0_11_add_566_6_lut (.I0(GND_net), .I1(n838[3]), 
            .I2(n604), .I3(n17179), .O(n837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_8 (.CI(n17058), .I0(n834[5]), .I1(n592), 
            .CO(n17059));
    SB_CARRY add_1234_5 (.CI(n17086), .I0(n835[14]), .I1(n747), .CO(n17087));
    SB_CARRY Alpha_15__I_0_11_add_566_6 (.CI(n17179), .I0(n838[3]), .I1(n604), 
            .CO(n17180));
    SB_LUT4 Alpha_15__I_0_11_add_566_5_lut (.I0(GND_net), .I1(n838[2]), 
            .I2(n604), .I3(n17178), .O(n837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_5 (.CI(n17178), .I0(n838[2]), .I1(n604), 
            .CO(n17179));
    SB_LUT4 Beta_15__I_0_add_562_7_lut (.I0(GND_net), .I1(n834[4]), .I2(n592), 
            .I3(n17057), .O(n833[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_566_4_lut (.I0(GND_net), .I1(n838[1]), 
            .I2(n604), .I3(n17177), .O(n837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_4 (.CI(n17177), .I0(n838[1]), .I1(n604), 
            .CO(n17178));
    SB_LUT4 Alpha_15__I_0_11_add_566_3_lut (.I0(GND_net), .I1(n838[0]), 
            .I2(n604), .I3(n17176), .O(n837[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_4_lut (.I0(GND_net), .I1(n834_adj_2173[14]), .I2(n743), 
            .I3(n17085), .O(Product1_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1234_4 (.CI(n17085), .I0(n834_adj_2173[14]), .I1(n743), 
            .CO(n17086));
    SB_CARRY Alpha_15__I_0_11_add_566_3 (.CI(n17176), .I0(n838[0]), .I1(n604), 
            .CO(n17177));
    SB_CARRY Beta_15__I_0_add_565_7 (.CI(n17012), .I0(n837_adj_2171[4]), 
            .I1(n601), .CO(n17013));
    SB_LUT4 Alpha_15__I_0_11_add_566_2_lut (.I0(GND_net), .I1(n607), .I2(n604), 
            .I3(GND_net), .O(n837[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_2 (.CI(GND_net), .I0(n607), .I1(n604), 
            .CO(n17176));
    SB_CARRY Beta_15__I_0_add_562_7 (.CI(n17057), .I0(n834[4]), .I1(n592), 
            .CO(n17058));
    SB_LUT4 Beta_15__I_0_add_564_12_lut (.I0(GND_net), .I1(n836[9]), .I2(n598), 
            .I3(n17032), .O(n835_adj_2172[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_14_lut (.I0(GND_net), .I1(n842[9]), .I2(n773), 
            .I3(n16946), .O(n841[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1232_2_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_out1_1[15]), 
            .I3(n16900), .O(Product4_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_2 (.CI(n16900), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[15]), 
            .CO(n16901));
    SB_LUT4 i11560_3_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(Look_Up_Table_out1_1[13]), .I3(GND_net), .O(n845[0]));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i11560_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 Alpha_15__I_0_11_i28_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n628));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Beta_15__I_0_i534_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n785));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i534_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Alpha_15__I_0_11_add_567_16_lut (.I0(GND_net), .I1(n839_adj_2174[13]), 
            .I2(n761), .I3(n17174), .O(n838[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_16 (.CI(n17174), .I0(n839_adj_2174[13]), 
            .I1(n761), .CO(n763));
    SB_LUT4 add_1234_3_lut (.I0(GND_net), .I1(n833_adj_2175[14]), .I2(n739), 
            .I3(n17084), .O(Product1_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_12 (.CI(n17032), .I0(n836[9]), .I1(n598), 
            .CO(n17033));
    SB_CARRY add_1234_3 (.CI(n17084), .I0(n833_adj_2175[14]), .I1(n739), 
            .CO(n17085));
    SB_LUT4 Beta_15__I_0_add_564_11_lut (.I0(GND_net), .I1(n836[8]), .I2(n598), 
            .I3(n17031), .O(n835_adj_2172[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_15_lut (.I0(GND_net), .I1(n841[11]), .I2(n613), 
            .I3(n16960), .O(n840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_11 (.CI(n17031), .I0(n836[8]), .I1(n598), 
            .CO(n17032));
    SB_LUT4 Beta_15__I_0_add_564_10_lut (.I0(GND_net), .I1(n836[7]), .I2(n598), 
            .I3(n17030), .O(n835_adj_2172[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_15 (.CI(n16960), .I0(n841[11]), .I1(n613), 
            .CO(n16961));
    SB_CARRY Beta_15__I_0_add_564_10 (.CI(n17030), .I0(n836[7]), .I1(n598), 
            .CO(n17031));
    SB_CARRY Beta_15__I_0_add_568_12 (.CI(n16972), .I0(n840[9]), .I1(n610), 
            .CO(n16973));
    SB_LUT4 Alpha_15__I_0_11_add_567_15_lut (.I0(GND_net), .I1(n839_adj_2174[12]), 
            .I2(n607), .I3(n17173), .O(n838[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_11_lut (.I0(GND_net), .I1(n839[8]), .I2(n607), 
            .I3(n16986), .O(n838_adj_2170[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_566_9_lut (.I0(GND_net), .I1(n838_adj_2170[6]), 
            .I2(n604), .I3(n16999), .O(n837_adj_2171[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_9_lut (.I0(GND_net), .I1(n836[6]), .I2(n598), 
            .I3(n17029), .O(n835_adj_2172[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_9 (.CI(n16999), .I0(n838_adj_2170[6]), 
            .I1(n604), .CO(n17000));
    SB_LUT4 Alpha_15__I_0_11_i10_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n601));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Beta_15__I_0_add_564_9 (.CI(n17029), .I0(n836[6]), .I1(n598), 
            .CO(n17030));
    SB_LUT4 Beta_15__I_0_add_564_8_lut (.I0(GND_net), .I1(n836[5]), .I2(n598), 
            .I3(n17028), .O(n835_adj_2172[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_15 (.CI(n17173), .I0(n839_adj_2174[12]), 
            .I1(n607), .CO(n17174));
    SB_CARRY Beta_15__I_0_add_564_8 (.CI(n17028), .I0(n836[5]), .I1(n598), 
            .CO(n17029));
    SB_LUT4 Beta_15__I_0_add_565_6_lut (.I0(GND_net), .I1(n837_adj_2171[3]), 
            .I2(n601), .I3(n17011), .O(n836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_7_lut (.I0(GND_net), .I1(n836[4]), .I2(n598), 
            .I3(n17027), .O(n835_adj_2172[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_2_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_out1_1[15]), 
            .I3(n17083), .O(Product1_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_6_lut (.I0(GND_net), .I1(n834[3]), .I2(n592), 
            .I3(n17056), .O(n833[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_567_14_lut (.I0(GND_net), .I1(n839_adj_2174[11]), 
            .I2(n607), .I3(n17172), .O(n838[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_7 (.CI(n17027), .I0(n836[4]), .I1(n598), 
            .CO(n17028));
    SB_LUT4 Beta_15__I_0_add_564_6_lut (.I0(GND_net), .I1(n836[3]), .I2(n598), 
            .I3(n17026), .O(n835_adj_2172[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_6 (.CI(n17056), .I0(n834[3]), .I1(n592), 
            .CO(n17057));
    SB_CARRY Alpha_15__I_0_11_add_567_14 (.CI(n17172), .I0(n839_adj_2174[11]), 
            .I1(n607), .CO(n17173));
    SB_LUT4 Alpha_15__I_0_11_add_567_13_lut (.I0(GND_net), .I1(n839_adj_2174[10]), 
            .I2(n607), .I3(n17171), .O(n838[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_11 (.CI(n16932), .I0(n843[7]), .I1(n619), 
            .CO(n16933));
    SB_CARRY Alpha_15__I_0_11_add_567_13 (.CI(n17171), .I0(n839_adj_2174[10]), 
            .I1(n607), .CO(n17172));
    SB_CARRY add_1234_2 (.CI(n17083), .I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[15]), 
            .CO(n17084));
    SB_LUT4 Alpha_15__I_0_11_add_567_12_lut (.I0(GND_net), .I1(n839_adj_2174[9]), 
            .I2(n607), .I3(n17170), .O(n838[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_12 (.CI(n17170), .I0(n839_adj_2174[9]), 
            .I1(n607), .CO(n17171));
    SB_CARRY add_1234_1 (.CI(GND_net), .I0(n832[14]), .I1(n832[14]), .CO(n17083));
    SB_LUT4 Beta_15__I_0_add_562_5_lut (.I0(GND_net), .I1(n834[2]), .I2(n592), 
            .I3(n17055), .O(n833[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_5 (.CI(n17055), .I0(n834[2]), .I1(n592), 
            .CO(n17056));
    SB_LUT4 Beta_15__I_0_add_561_16_lut (.I0(GND_net), .I1(n833[13]), .I2(n737), 
            .I3(n17081), .O(n832_adj_2176[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_567_11_lut (.I0(GND_net), .I1(n839_adj_2174[8]), 
            .I2(n607), .I3(n17169), .O(n838[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_16 (.CI(n17081), .I0(n833[13]), .I1(n737), 
            .CO(n739_adj_2006));
    SB_CARRY Beta_15__I_0_add_564_6 (.CI(n17026), .I0(n836[3]), .I1(n598), 
            .CO(n17027));
    SB_LUT4 Beta_15__I_0_add_562_4_lut (.I0(GND_net), .I1(n834[1]), .I2(n592), 
            .I3(n17054), .O(n833[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1232_13_lut (.I0(GND_net), .I1(n843[14]), .I2(n779), .I3(n16911), 
            .O(Product4_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_4 (.CI(n17054), .I0(n834[1]), .I1(n592), 
            .CO(n17055));
    SB_LUT4 Beta_15__I_0_add_568_11_lut (.I0(GND_net), .I1(n840[8]), .I2(n610), 
            .I3(n16971), .O(n839[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_11 (.CI(n16986), .I0(n839[8]), .I1(n607), 
            .CO(n16987));
    SB_LUT4 Beta_15__I_0_add_567_10_lut (.I0(GND_net), .I1(n839[7]), .I2(n607), 
            .I3(n16985), .O(n838_adj_2170[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_3_lut (.I0(GND_net), .I1(n834[0]), .I2(n592), 
            .I3(n17053), .O(n833[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_11 (.CI(n17169), .I0(n839_adj_2174[8]), 
            .I1(n607), .CO(n17170));
    SB_LUT4 Alpha_15__I_0_11_add_567_10_lut (.I0(GND_net), .I1(n839_adj_2174[7]), 
            .I2(n607), .I3(n17168), .O(n838[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_3 (.CI(n17053), .I0(n834[0]), .I1(n592), 
            .CO(n17054));
    SB_LUT4 Beta_15__I_0_add_566_8_lut (.I0(GND_net), .I1(n838_adj_2170[5]), 
            .I2(n604), .I3(n16998), .O(n837_adj_2171[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_10 (.CI(n17168), .I0(n839_adj_2174[7]), 
            .I1(n607), .CO(n17169));
    SB_CARRY Beta_15__I_0_add_565_6 (.CI(n17011), .I0(n837_adj_2171[3]), 
            .I1(n601), .CO(n17012));
    SB_LUT4 Alpha_15__I_0_11_add_567_9_lut (.I0(GND_net), .I1(n839_adj_2174[6]), 
            .I2(n607), .I3(n17167), .O(n838[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_5_lut (.I0(GND_net), .I1(n836[2]), .I2(n598), 
            .I3(n17025), .O(n835_adj_2172[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_5 (.CI(n17025), .I0(n836[2]), .I1(n598), 
            .CO(n17026));
    SB_LUT4 Beta_15__I_0_add_561_15_lut (.I0(GND_net), .I1(n833[12]), .I2(dCurrent[2]), 
            .I3(n17080), .O(Product4_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_2_lut (.I0(GND_net), .I1(n595), .I2(n592), 
            .I3(GND_net), .O(n833[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_15 (.CI(n17080), .I0(n833[12]), .I1(dCurrent[2]), 
            .CO(n17081));
    SB_LUT4 Beta_15__I_0_add_564_4_lut (.I0(GND_net), .I1(n836[1]), .I2(n598), 
            .I3(n17024), .O(n835_adj_2172[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_9 (.CI(n17167), .I0(n839_adj_2174[6]), 
            .I1(n607), .CO(n17168));
    SB_LUT4 Beta_15__I_0_add_561_14_lut (.I0(GND_net), .I1(n833[11]), .I2(dCurrent[2]), 
            .I3(n17079), .O(Product4_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_567_8_lut (.I0(GND_net), .I1(n839_adj_2174[5]), 
            .I2(n607), .I3(n17166), .O(n838[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_2 (.CI(GND_net), .I0(n595), .I1(n592), 
            .CO(n17053));
    SB_LUT4 Beta_15__I_0_add_569_14_lut (.I0(GND_net), .I1(n841[11]), .I2(n613), 
            .I3(n16959), .O(n840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_563_16_lut (.I0(GND_net), .I1(n835_adj_2172[13]), 
            .I2(n745), .I3(n17051), .O(n834[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_16 (.CI(n17051), .I0(n835_adj_2172[13]), 
            .I1(n745), .CO(n747_adj_2012));
    SB_LUT4 Beta_15__I_0_add_572_9_lut (.I0(GND_net), .I1(n844[5]), .I2(n622), 
            .I3(n16921), .O(n843[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_8 (.CI(n17166), .I0(n839_adj_2174[5]), 
            .I1(n607), .CO(n17167));
    SB_LUT4 Alpha_15__I_0_11_add_567_7_lut (.I0(GND_net), .I1(n839_adj_2174[4]), 
            .I2(n607), .I3(n17165), .O(n838[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_563_15_lut (.I0(GND_net), .I1(n835_adj_2172[12]), 
            .I2(n595), .I3(n17050), .O(n834[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_10_lut (.I0(GND_net), .I1(n843[7]), .I2(n619), 
            .I3(n16931), .O(n842[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_15 (.CI(n17050), .I0(n835_adj_2172[12]), 
            .I1(n595), .CO(n17051));
    SB_CARRY Beta_15__I_0_add_561_14 (.CI(n17079), .I0(n833[11]), .I1(dCurrent[2]), 
            .CO(n17080));
    SB_LUT4 Beta_15__I_0_add_561_13_lut (.I0(GND_net), .I1(n833[10]), .I2(dCurrent[2]), 
            .I3(n17078), .O(Product4_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_7 (.CI(n17165), .I0(n839_adj_2174[4]), 
            .I1(n607), .CO(n17166));
    SB_LUT4 Alpha_15__I_0_11_add_567_6_lut (.I0(GND_net), .I1(n839_adj_2174[3]), 
            .I2(n607), .I3(n17164), .O(n838[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_6 (.CI(n17164), .I0(n839_adj_2174[3]), 
            .I1(n607), .CO(n17165));
    SB_CARRY Beta_15__I_0_add_572_9 (.CI(n16921), .I0(n844[5]), .I1(n622), 
            .CO(n16922));
    SB_LUT4 Alpha_15__I_0_11_add_567_5_lut (.I0(GND_net), .I1(n839_adj_2174[2]), 
            .I2(n607), .I3(n17163), .O(n838[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_1 (.CI(GND_net), .I0(n832_adj_2176[14]), .I1(n832_adj_2176[14]), 
            .CO(n16900));
    SB_CARRY add_1232_13 (.CI(n16911), .I0(n843[14]), .I1(n779), .CO(n16912));
    SB_LUT4 add_1232_12_lut (.I0(GND_net), .I1(n842[14]), .I2(n775), .I3(n16910), 
            .O(Product4_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_5 (.CI(n17163), .I0(n839_adj_2174[2]), 
            .I1(n607), .CO(n17164));
    SB_LUT4 Beta_15__I_0_add_572_8_lut (.I0(GND_net), .I1(n844[5]), .I2(n622), 
            .I3(n16920), .O(n843[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_10 (.CI(n16931), .I0(n843[7]), .I1(n619), 
            .CO(n16932));
    SB_CARRY Beta_15__I_0_add_570_14 (.CI(n16946), .I0(n842[9]), .I1(n773), 
            .CO(n775));
    SB_LUT4 Beta_15__I_0_add_571_9_lut (.I0(GND_net), .I1(n843[6]), .I2(n619), 
            .I3(n16930), .O(n842[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_13_lut (.I0(GND_net), .I1(n842[9]), .I2(n616), 
            .I3(n16945), .O(n841[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_567_4_lut (.I0(GND_net), .I1(n839_adj_2174[1]), 
            .I2(n607), .I3(n17162), .O(n838[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_14 (.CI(n16959), .I0(n841[11]), .I1(n613), 
            .CO(n16960));
    SB_CARRY Beta_15__I_0_add_568_11 (.CI(n16971), .I0(n840[8]), .I1(n610), 
            .CO(n16972));
    SB_CARRY Beta_15__I_0_add_567_10 (.CI(n16985), .I0(n839[7]), .I1(n607), 
            .CO(n16986));
    SB_LUT4 Beta_15__I_0_add_567_9_lut (.I0(GND_net), .I1(n839[6]), .I2(n607), 
            .I3(n16984), .O(n838_adj_2170[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_4 (.CI(n17162), .I0(n839_adj_2174[1]), 
            .I1(n607), .CO(n17163));
    SB_CARRY Beta_15__I_0_add_566_8 (.CI(n16998), .I0(n838_adj_2170[5]), 
            .I1(n604), .CO(n16999));
    SB_LUT4 Beta_15__I_0_add_565_5_lut (.I0(GND_net), .I1(n837_adj_2171[2]), 
            .I2(n601), .I3(n17010), .O(n836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_4 (.CI(n17024), .I0(n836[1]), .I1(n598), 
            .CO(n17025));
    SB_LUT4 Beta_15__I_0_add_564_3_lut (.I0(GND_net), .I1(n836[0]), .I2(n598), 
            .I3(n17023), .O(n835_adj_2172[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_9 (.CI(n16930), .I0(n843[6]), .I1(n619), 
            .CO(n16931));
    SB_CARRY Beta_15__I_0_add_570_13 (.CI(n16945), .I0(n842[9]), .I1(n616), 
            .CO(n16946));
    SB_LUT4 Alpha_15__I_0_11_add_567_3_lut (.I0(GND_net), .I1(n839_adj_2174[0]), 
            .I2(n607), .I3(n17161), .O(n838[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_563_14_lut (.I0(GND_net), .I1(n835_adj_2172[11]), 
            .I2(n595), .I3(n17049), .O(n834[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_13 (.CI(n17078), .I0(n833[10]), .I1(dCurrent[2]), 
            .CO(n17079));
    SB_CARRY Alpha_15__I_0_11_add_567_3 (.CI(n17161), .I0(n839_adj_2174[0]), 
            .I1(n607), .CO(n17162));
    SB_LUT4 Alpha_15__I_0_11_add_567_2_lut (.I0(GND_net), .I1(n610), .I2(n607), 
            .I3(GND_net), .O(n838[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_567_2 (.CI(GND_net), .I0(n610), .I1(n607), 
            .CO(n17161));
    SB_LUT4 Alpha_15__I_0_11_add_568_16_lut (.I0(GND_net), .I1(n840_adj_2177[13]), 
            .I2(n765), .I3(n17159), .O(n839_adj_2174[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_16 (.CI(n17159), .I0(n840_adj_2177[13]), 
            .I1(n765), .CO(n767));
    SB_LUT4 Beta_15__I_0_add_569_13_lut (.I0(GND_net), .I1(n841[10]), .I2(n613), 
            .I3(n16958), .O(n840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_14 (.CI(n17049), .I0(n835_adj_2172[11]), 
            .I1(n595), .CO(n17050));
    SB_LUT4 Beta_15__I_0_add_571_8_lut (.I0(GND_net), .I1(n843[5]), .I2(n619), 
            .I3(n16929), .O(n842[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_13 (.CI(n16958), .I0(n841[10]), .I1(n613), 
            .CO(n16959));
    SB_LUT4 Alpha_15__I_0_11_add_568_15_lut (.I0(GND_net), .I1(n840_adj_2177[12]), 
            .I2(n610), .I3(n17158), .O(n839_adj_2174[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_15 (.CI(n17158), .I0(n840_adj_2177[12]), 
            .I1(n610), .CO(n17159));
    SB_LUT4 Alpha_15__I_0_11_add_568_14_lut (.I0(GND_net), .I1(n840_adj_2177[11]), 
            .I2(n610), .I3(n17157), .O(n839_adj_2174[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_14 (.CI(n17157), .I0(n840_adj_2177[11]), 
            .I1(n610), .CO(n17158));
    SB_LUT4 Alpha_15__I_0_11_add_568_13_lut (.I0(GND_net), .I1(n840_adj_2177[10]), 
            .I2(n610), .I3(n17156), .O(n839_adj_2174[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_13 (.CI(n17156), .I0(n840_adj_2177[10]), 
            .I1(n610), .CO(n17157));
    SB_CARRY add_1232_12 (.CI(n16910), .I0(n842[14]), .I1(n775), .CO(n16911));
    SB_LUT4 add_1232_11_lut (.I0(GND_net), .I1(n841[14]), .I2(n771), .I3(n16909), 
            .O(Product4_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_568_12_lut (.I0(GND_net), .I1(n840_adj_2177[9]), 
            .I2(n610), .I3(n17155), .O(n839_adj_2174[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_8 (.CI(n16920), .I0(n844[5]), .I1(n622), 
            .CO(n16921));
    SB_LUT4 Beta_15__I_0_add_570_12_lut (.I0(GND_net), .I1(n842[9]), .I2(n616), 
            .I3(n16944), .O(n841[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_12 (.CI(n16944), .I0(n842[9]), .I1(n616), 
            .CO(n16945));
    SB_CARRY Alpha_15__I_0_11_add_568_12 (.CI(n17155), .I0(n840_adj_2177[9]), 
            .I1(n610), .CO(n17156));
    SB_LUT4 Alpha_15__I_0_11_add_568_11_lut (.I0(GND_net), .I1(n840_adj_2177[8]), 
            .I2(n610), .I3(n17154), .O(n839_adj_2174[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_10_lut (.I0(GND_net), .I1(n840[7]), .I2(n610), 
            .I3(n16970), .O(n839[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_12_lut (.I0(GND_net), .I1(n841[9]), .I2(n613), 
            .I3(n16957), .O(n840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_10 (.CI(n16970), .I0(n840[7]), .I1(n610), 
            .CO(n16971));
    SB_CARRY Beta_15__I_0_add_567_9 (.CI(n16984), .I0(n839[6]), .I1(n607), 
            .CO(n16985));
    SB_LUT4 Beta_15__I_0_add_567_8_lut (.I0(GND_net), .I1(n839[5]), .I2(n607), 
            .I3(n16983), .O(n838_adj_2170[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_11 (.CI(n17154), .I0(n840_adj_2177[8]), 
            .I1(n610), .CO(n17155));
    SB_LUT4 Beta_15__I_0_add_566_7_lut (.I0(GND_net), .I1(n838_adj_2170[4]), 
            .I2(n604), .I3(n16997), .O(n837_adj_2171[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_5 (.CI(n17010), .I0(n837_adj_2171[2]), 
            .I1(n601), .CO(n17011));
    SB_CARRY Beta_15__I_0_add_564_3 (.CI(n17023), .I0(n836[0]), .I1(n598), 
            .CO(n17024));
    SB_CARRY Beta_15__I_0_add_571_8 (.CI(n16929), .I0(n843[5]), .I1(n619), 
            .CO(n16930));
    SB_LUT4 Alpha_15__I_0_11_add_568_10_lut (.I0(GND_net), .I1(n840_adj_2177[7]), 
            .I2(n610), .I3(n17153), .O(n839_adj_2174[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_563_13_lut (.I0(GND_net), .I1(n835_adj_2172[10]), 
            .I2(n595), .I3(n17048), .O(n834[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_8 (.CI(n16983), .I0(n839[5]), .I1(n607), 
            .CO(n16984));
    SB_LUT4 Beta_15__I_0_add_561_12_lut (.I0(GND_net), .I1(n833[9]), .I2(dCurrent[2]), 
            .I3(n17077), .O(Product4_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_10 (.CI(n17153), .I0(n840_adj_2177[7]), 
            .I1(n610), .CO(n17154));
    SB_LUT4 Alpha_15__I_0_11_add_568_9_lut (.I0(GND_net), .I1(n840_adj_2177[6]), 
            .I2(n610), .I3(n17152), .O(n839_adj_2174[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_9 (.CI(n17152), .I0(n840_adj_2177[6]), 
            .I1(n610), .CO(n17153));
    SB_CARRY Beta_15__I_0_add_566_7 (.CI(n16997), .I0(n838_adj_2170[4]), 
            .I1(n604), .CO(n16998));
    SB_CARRY Beta_15__I_0_add_561_12 (.CI(n17077), .I0(n833[9]), .I1(dCurrent[2]), 
            .CO(n17078));
    SB_LUT4 Beta_15__I_0_add_566_6_lut (.I0(GND_net), .I1(n838_adj_2170[3]), 
            .I2(n604), .I3(n16996), .O(n837_adj_2171[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_568_8_lut (.I0(GND_net), .I1(n840_adj_2177[5]), 
            .I2(n610), .I3(n17151), .O(n839_adj_2174[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_8 (.CI(n17151), .I0(n840_adj_2177[5]), 
            .I1(n610), .CO(n17152));
    SB_LUT4 Alpha_15__I_0_11_add_568_7_lut (.I0(GND_net), .I1(n840_adj_2177[4]), 
            .I2(n610), .I3(n17150), .O(n839_adj_2174[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_7 (.CI(n17150), .I0(n840_adj_2177[4]), 
            .I1(n610), .CO(n17151));
    SB_LUT4 Alpha_15__I_0_11_add_568_6_lut (.I0(GND_net), .I1(n840_adj_2177[3]), 
            .I2(n610), .I3(n17149), .O(n839_adj_2174[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_561_11_lut (.I0(GND_net), .I1(n833[8]), .I2(dCurrent[2]), 
            .I3(n17076), .O(Product4_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_11 (.CI(n16909), .I0(n841[14]), .I1(n771), .CO(n16910));
    SB_LUT4 Beta_15__I_0_add_572_7_lut (.I0(GND_net), .I1(n844[4]), .I2(n622), 
            .I3(n16919), .O(n843[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_7 (.CI(n16919), .I0(n844[4]), .I1(n622), 
            .CO(n16920));
    SB_CARRY Alpha_15__I_0_11_add_568_6 (.CI(n17149), .I0(n840_adj_2177[3]), 
            .I1(n610), .CO(n17150));
    SB_LUT4 Beta_15__I_0_add_571_7_lut (.I0(GND_net), .I1(n843[4]), .I2(n619), 
            .I3(n16928), .O(n842[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_11_lut (.I0(GND_net), .I1(n842[8]), .I2(n616), 
            .I3(n16943), .O(n841[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_12 (.CI(n16957), .I0(n841[9]), .I1(n613), 
            .CO(n16958));
    SB_LUT4 Beta_15__I_0_add_569_11_lut (.I0(GND_net), .I1(n841[8]), .I2(n613), 
            .I3(n16956), .O(n840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_568_5_lut (.I0(GND_net), .I1(n840_adj_2177[2]), 
            .I2(n610), .I3(n17148), .O(n839_adj_2174[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_9_lut (.I0(GND_net), .I1(n840[6]), .I2(n610), 
            .I3(n16969), .O(n839[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_7_lut (.I0(GND_net), .I1(n839[4]), .I2(n607), 
            .I3(n16982), .O(n838_adj_2170[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_5 (.CI(n17148), .I0(n840_adj_2177[2]), 
            .I1(n610), .CO(n17149));
    SB_LUT4 Beta_15__I_0_add_564_2_lut (.I0(GND_net), .I1(n601), .I2(n598), 
            .I3(GND_net), .O(n835_adj_2172[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_565_4_lut (.I0(GND_net), .I1(n837_adj_2171[1]), 
            .I2(n601), .I3(n17009), .O(n836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_568_4_lut (.I0(GND_net), .I1(n840_adj_2177[1]), 
            .I2(n610), .I3(n17147), .O(n839_adj_2174[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_4 (.CI(n17147), .I0(n840_adj_2177[1]), 
            .I1(n610), .CO(n17148));
    SB_CARRY Beta_15__I_0_add_563_13 (.CI(n17048), .I0(n835_adj_2172[10]), 
            .I1(n595), .CO(n17049));
    SB_LUT4 Beta_15__I_0_add_563_12_lut (.I0(GND_net), .I1(n835_adj_2172[9]), 
            .I2(n595), .I3(n17047), .O(n834[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_12 (.CI(n17047), .I0(n835_adj_2172[9]), 
            .I1(n595), .CO(n17048));
    SB_LUT4 Beta_15__I_0_add_563_11_lut (.I0(GND_net), .I1(n835_adj_2172[8]), 
            .I2(n595), .I3(n17046), .O(n834[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_11 (.CI(n17046), .I0(n835_adj_2172[8]), 
            .I1(n595), .CO(n17047));
    SB_LUT4 Beta_15__I_0_add_563_10_lut (.I0(GND_net), .I1(n835_adj_2172[7]), 
            .I2(n595), .I3(n17045), .O(n834[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_10 (.CI(n17045), .I0(n835_adj_2172[7]), 
            .I1(n595), .CO(n17046));
    SB_LUT4 Alpha_15__I_0_11_add_568_3_lut (.I0(GND_net), .I1(n840_adj_2177[0]), 
            .I2(n610), .I3(n17146), .O(n839_adj_2174[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_3 (.CI(n17146), .I0(n840_adj_2177[0]), 
            .I1(n610), .CO(n17147));
    SB_LUT4 Beta_15__I_0_add_563_9_lut (.I0(GND_net), .I1(n835_adj_2172[6]), 
            .I2(n595), .I3(n17044), .O(n834[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_11 (.CI(n17076), .I0(n833[8]), .I1(dCurrent[2]), 
            .CO(n17077));
    SB_CARRY Beta_15__I_0_add_566_6 (.CI(n16996), .I0(n838_adj_2170[3]), 
            .I1(n604), .CO(n16997));
    SB_LUT4 Beta_15__I_0_add_566_5_lut (.I0(GND_net), .I1(n838_adj_2170[2]), 
            .I2(n604), .I3(n16995), .O(n837_adj_2171[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_9 (.CI(n17044), .I0(n835_adj_2172[6]), 
            .I1(n595), .CO(n17045));
    SB_LUT4 Alpha_15__I_0_11_add_568_2_lut (.I0(GND_net), .I1(n613), .I2(n610), 
            .I3(GND_net), .O(n839_adj_2174[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_568_2 (.CI(GND_net), .I0(n613), .I1(n610), 
            .CO(n17146));
    SB_LUT4 Alpha_15__I_0_11_add_569_16_lut (.I0(GND_net), .I1(n841_adj_2178[11]), 
            .I2(n769), .I3(n17144), .O(n840_adj_2177[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_4 (.CI(n17009), .I0(n837_adj_2171[1]), 
            .I1(n601), .CO(n17010));
    SB_CARRY Alpha_15__I_0_11_add_569_16 (.CI(n17144), .I0(n841_adj_2178[11]), 
            .I1(n769), .CO(n771_adj_2032));
    SB_LUT4 Beta_15__I_0_add_561_10_lut (.I0(GND_net), .I1(n833[7]), .I2(dCurrent[2]), 
            .I3(n17075), .O(Product4_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_2 (.CI(GND_net), .I0(n601), .I1(n598), 
            .CO(n17023));
    SB_LUT4 Alpha_15__I_0_11_add_569_15_lut (.I0(GND_net), .I1(n841_adj_2178[11]), 
            .I2(n613), .I3(n17143), .O(n840_adj_2177[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_11 (.CI(n16956), .I0(n841[8]), .I1(n613), 
            .CO(n16957));
    SB_CARRY Alpha_15__I_0_11_add_569_15 (.CI(n17143), .I0(n841_adj_2178[11]), 
            .I1(n613), .CO(n17144));
    SB_LUT4 Beta_15__I_0_add_563_8_lut (.I0(GND_net), .I1(n835_adj_2172[5]), 
            .I2(n595), .I3(n17043), .O(n834[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_569_14_lut (.I0(GND_net), .I1(n841_adj_2178[11]), 
            .I2(n613), .I3(n17142), .O(n840_adj_2177[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_8 (.CI(n17043), .I0(n835_adj_2172[5]), 
            .I1(n595), .CO(n17044));
    SB_LUT4 Beta_15__I_0_add_569_10_lut (.I0(GND_net), .I1(n841[7]), .I2(n613), 
            .I3(n16955), .O(n840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_9 (.CI(n16969), .I0(n840[6]), .I1(n610), 
            .CO(n16970));
    SB_CARRY Beta_15__I_0_add_567_7 (.CI(n16982), .I0(n839[4]), .I1(n607), 
            .CO(n16983));
    SB_LUT4 Beta_15__I_0_add_565_3_lut (.I0(GND_net), .I1(n837_adj_2171[0]), 
            .I2(n601), .I3(n17008), .O(n836[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_14 (.CI(n17142), .I0(n841_adj_2178[11]), 
            .I1(n613), .CO(n17143));
    SB_CARRY Beta_15__I_0_add_561_10 (.CI(n17075), .I0(n833[7]), .I1(dCurrent[2]), 
            .CO(n17076));
    SB_LUT4 Beta_15__I_0_add_561_9_lut (.I0(GND_net), .I1(n833[6]), .I2(dCurrent[2]), 
            .I3(n17074), .O(Product4_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_3 (.CI(n17008), .I0(n837_adj_2171[0]), 
            .I1(n601), .CO(n17009));
    SB_LUT4 Alpha_15__I_0_11_add_569_13_lut (.I0(GND_net), .I1(n841_adj_2178[10]), 
            .I2(n613), .I3(n17141), .O(n840_adj_2177[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_9 (.CI(n17074), .I0(n833[6]), .I1(dCurrent[2]), 
            .CO(n17075));
    SB_CARRY Alpha_15__I_0_11_add_569_13 (.CI(n17141), .I0(n841_adj_2178[10]), 
            .I1(n613), .CO(n17142));
    SB_CARRY Beta_15__I_0_add_570_11 (.CI(n16943), .I0(n842[8]), .I1(n616), 
            .CO(n16944));
    SB_LUT4 Beta_15__I_0_add_561_8_lut (.I0(GND_net), .I1(n833[5]), .I2(dCurrent[2]), 
            .I3(n17073), .O(Product4_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_8 (.CI(n17073), .I0(n833[5]), .I1(dCurrent[2]), 
            .CO(n17074));
    SB_LUT4 Beta_15__I_0_add_570_10_lut (.I0(GND_net), .I1(n842[7]), .I2(n616), 
            .I3(n16942), .O(n841[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_565_16_lut (.I0(GND_net), .I1(n837_adj_2171[13]), 
            .I2(n753), .I3(n17021), .O(n836[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_569_12_lut (.I0(GND_net), .I1(n841_adj_2178[9]), 
            .I2(n613), .I3(n17140), .O(n840_adj_2177[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_561_7_lut (.I0(GND_net), .I1(n833[4]), .I2(dCurrent[2]), 
            .I3(n17072), .O(Product4_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_5 (.CI(n16995), .I0(n838_adj_2170[2]), 
            .I1(n604), .CO(n16996));
    SB_LUT4 Beta_15__I_0_add_568_8_lut (.I0(GND_net), .I1(n840[5]), .I2(n610), 
            .I3(n16968), .O(n839[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_12 (.CI(n17140), .I0(n841_adj_2178[9]), 
            .I1(n613), .CO(n17141));
    SB_LUT4 Beta_15__I_0_add_566_4_lut (.I0(GND_net), .I1(n838_adj_2170[1]), 
            .I2(n604), .I3(n16994), .O(n837_adj_2171[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_569_11_lut (.I0(GND_net), .I1(n841_adj_2178[8]), 
            .I2(n613), .I3(n17139), .O(n840_adj_2177[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_11 (.CI(n17139), .I0(n841_adj_2178[8]), 
            .I1(n613), .CO(n17140));
    SB_LUT4 Beta_15__I_0_add_565_2_lut (.I0(GND_net), .I1(n604), .I2(n601), 
            .I3(GND_net), .O(n836[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_7 (.CI(n17072), .I0(n833[4]), .I1(dCurrent[2]), 
            .CO(n17073));
    SB_LUT4 Alpha_15__I_0_11_add_569_10_lut (.I0(GND_net), .I1(n841_adj_2178[7]), 
            .I2(n613), .I3(n17138), .O(n840_adj_2177[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_10 (.CI(n17138), .I0(n841_adj_2178[7]), 
            .I1(n613), .CO(n17139));
    SB_CARRY Beta_15__I_0_add_570_10 (.CI(n16942), .I0(n842[7]), .I1(n616), 
            .CO(n16943));
    SB_LUT4 Alpha_15__I_0_11_add_569_9_lut (.I0(GND_net), .I1(n841_adj_2178[6]), 
            .I2(n613), .I3(n17137), .O(n840_adj_2177[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_9 (.CI(n17137), .I0(n841_adj_2178[6]), 
            .I1(n613), .CO(n17138));
    SB_LUT4 Beta_15__I_0_add_567_6_lut (.I0(GND_net), .I1(n839[3]), .I2(n607), 
            .I3(n16981), .O(n838_adj_2170[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_9_lut (.I0(GND_net), .I1(n842[6]), .I2(n616), 
            .I3(n16941), .O(n841[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_569_8_lut (.I0(GND_net), .I1(n841_adj_2178[5]), 
            .I2(n613), .I3(n17136), .O(n840_adj_2177[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_8 (.CI(n17136), .I0(n841_adj_2178[5]), 
            .I1(n613), .CO(n17137));
    SB_LUT4 Alpha_15__I_0_11_add_569_7_lut (.I0(GND_net), .I1(n841_adj_2178[4]), 
            .I2(n613), .I3(n17135), .O(n840_adj_2177[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_7 (.CI(n17135), .I0(n841_adj_2178[4]), 
            .I1(n613), .CO(n17136));
    SB_LUT4 Alpha_15__I_0_11_add_569_6_lut (.I0(GND_net), .I1(n841_adj_2178[3]), 
            .I2(n613), .I3(n17134), .O(n840_adj_2177[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_10 (.CI(n16955), .I0(n841[7]), .I1(n613), 
            .CO(n16956));
    SB_CARRY Alpha_15__I_0_11_add_569_6 (.CI(n17134), .I0(n841_adj_2178[3]), 
            .I1(n613), .CO(n17135));
    SB_LUT4 Alpha_15__I_0_11_add_569_5_lut (.I0(GND_net), .I1(n841_adj_2178[2]), 
            .I2(n613), .I3(n17133), .O(n840_adj_2177[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_5 (.CI(n17133), .I0(n841_adj_2178[2]), 
            .I1(n613), .CO(n17134));
    SB_LUT4 add_1232_10_lut (.I0(GND_net), .I1(n840[14]), .I2(n767_adj_2041), 
            .I3(n16908), .O(Product4_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_572_6_lut (.I0(GND_net), .I1(n844[3]), .I2(n622), 
            .I3(n16918), .O(n843[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_7 (.CI(n16928), .I0(n843[4]), .I1(n619), 
            .CO(n16929));
    SB_LUT4 Alpha_15__I_0_11_add_569_4_lut (.I0(GND_net), .I1(n841_adj_2178[1]), 
            .I2(n613), .I3(n17132), .O(n840_adj_2177[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_6_lut (.I0(GND_net), .I1(n843[3]), .I2(n619), 
            .I3(n16927), .O(n842[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_4 (.CI(n17132), .I0(n841_adj_2178[1]), 
            .I1(n613), .CO(n17133));
    SB_CARRY Beta_15__I_0_add_570_9 (.CI(n16941), .I0(n842[6]), .I1(n616), 
            .CO(n16942));
    SB_LUT4 Beta_15__I_0_add_569_9_lut (.I0(GND_net), .I1(n841[6]), .I2(n613), 
            .I3(n16954), .O(n840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_8 (.CI(n16968), .I0(n840[5]), .I1(n610), 
            .CO(n16969));
    SB_LUT4 Beta_15__I_0_add_568_7_lut (.I0(GND_net), .I1(n840[4]), .I2(n610), 
            .I3(n16967), .O(n839[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_569_3_lut (.I0(GND_net), .I1(n841_adj_2178[0]), 
            .I2(n613), .I3(n17131), .O(n840_adj_2177[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_6 (.CI(n16981), .I0(n839[3]), .I1(n607), 
            .CO(n16982));
    SB_CARRY Beta_15__I_0_add_566_4 (.CI(n16994), .I0(n838_adj_2170[1]), 
            .I1(n604), .CO(n16995));
    SB_CARRY Beta_15__I_0_add_565_2 (.CI(GND_net), .I0(n604), .I1(n601), 
            .CO(n17008));
    SB_LUT4 Beta_15__I_0_add_566_16_lut (.I0(GND_net), .I1(n838_adj_2170[13]), 
            .I2(n757), .I3(n17006), .O(n837_adj_2171[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_3 (.CI(n17131), .I0(n841_adj_2178[0]), 
            .I1(n613), .CO(n17132));
    SB_CARRY Beta_15__I_0_add_565_16 (.CI(n17021), .I0(n837_adj_2171[13]), 
            .I1(n753), .CO(n755));
    SB_LUT4 Beta_15__I_0_add_563_7_lut (.I0(GND_net), .I1(n835_adj_2172[4]), 
            .I2(n595), .I3(n17042), .O(n834[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_7 (.CI(n17042), .I0(n835_adj_2172[4]), 
            .I1(n595), .CO(n17043));
    SB_LUT4 Beta_15__I_0_add_561_6_lut (.I0(GND_net), .I1(n833[3]), .I2(dCurrent[2]), 
            .I3(n17071), .O(Product4_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_569_2_lut (.I0(GND_net), .I1(n616), .I2(n613), 
            .I3(GND_net), .O(n840_adj_2177[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_569_2 (.CI(GND_net), .I0(n616), .I1(n613), 
            .CO(n17131));
    SB_LUT4 Alpha_15__I_0_11_add_570_14_lut (.I0(GND_net), .I1(n842_adj_2179[9]), 
            .I2(n773), .I3(n17129), .O(n841_adj_2178[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_6 (.CI(n17071), .I0(n833[3]), .I1(dCurrent[2]), 
            .CO(n17072));
    SB_CARRY Alpha_15__I_0_11_add_570_14 (.CI(n17129), .I0(n842_adj_2179[9]), 
            .I1(n773), .CO(n775_adj_2047));
    SB_LUT4 Beta_15__I_0_add_561_5_lut (.I0(GND_net), .I1(n833[2]), .I2(dCurrent[2]), 
            .I3(n17070), .O(Product4_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_7 (.CI(n16967), .I0(n840[4]), .I1(n610), 
            .CO(n16968));
    SB_LUT4 Beta_15__I_0_add_565_15_lut (.I0(GND_net), .I1(n837_adj_2171[12]), 
            .I2(n601), .I3(n17020), .O(n836[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_29_lut (.I0(GND_net), .I1(Product1_mul_temp[29]), .I2(GND_net), 
            .I3(n17303), .O(\dCurrent[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_28_lut (.I0(GND_net), .I1(Product1_mul_temp[28]), .I2(GND_net), 
            .I3(n17302), .O(\dCurrent[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_28 (.CI(n17302), .I0(Product1_mul_temp[28]), .I1(GND_net), 
            .CO(n17303));
    SB_LUT4 add_8094_27_lut (.I0(GND_net), .I1(Product1_mul_temp[27]), .I2(GND_net), 
            .I3(n17301), .O(\dCurrent[29] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_27 (.CI(n17301), .I0(Product1_mul_temp[27]), .I1(GND_net), 
            .CO(n17302));
    SB_LUT4 add_8094_26_lut (.I0(GND_net), .I1(Product1_mul_temp[26]), .I2(GND_net), 
            .I3(n17300), .O(\dCurrent[28] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_26 (.CI(n17300), .I0(Product1_mul_temp[26]), .I1(GND_net), 
            .CO(n17301));
    SB_LUT4 add_8094_25_lut (.I0(GND_net), .I1(Product1_mul_temp[25]), .I2(GND_net), 
            .I3(n17299), .O(\dCurrent[27] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_25 (.CI(n17299), .I0(Product1_mul_temp[25]), .I1(GND_net), 
            .CO(n17300));
    SB_LUT4 add_8094_24_lut (.I0(GND_net), .I1(Product1_mul_temp[24]), .I2(GND_net), 
            .I3(n17298), .O(\dCurrent[26] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_24 (.CI(n17298), .I0(Product1_mul_temp[24]), .I1(GND_net), 
            .CO(n17299));
    SB_LUT4 add_8094_23_lut (.I0(GND_net), .I1(Product1_mul_temp[23]), .I2(GND_net), 
            .I3(n17297), .O(\dCurrent[25] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_23 (.CI(n17297), .I0(Product1_mul_temp[23]), .I1(GND_net), 
            .CO(n17298));
    SB_LUT4 Alpha_15__I_0_11_add_570_13_lut (.I0(GND_net), .I1(n842_adj_2179[9]), 
            .I2(n616), .I3(n17128), .O(n841_adj_2178[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_22_lut (.I0(GND_net), .I1(Product1_mul_temp[22]), .I2(GND_net), 
            .I3(n17296), .O(\dCurrent[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_13 (.CI(n17128), .I0(n842_adj_2179[9]), 
            .I1(n616), .CO(n17129));
    SB_CARRY add_8094_22 (.CI(n17296), .I0(Product1_mul_temp[22]), .I1(GND_net), 
            .CO(n17297));
    SB_LUT4 Beta_15__I_0_add_567_5_lut (.I0(GND_net), .I1(n839[2]), .I2(n607), 
            .I3(n16980), .O(n838_adj_2170[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_8_lut (.I0(GND_net), .I1(n842[5]), .I2(n616), 
            .I3(n16940), .O(n841[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_21_lut (.I0(GND_net), .I1(Product1_mul_temp[21]), .I2(GND_net), 
            .I3(n17295), .O(\dCurrent[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_570_12_lut (.I0(GND_net), .I1(n842_adj_2179[9]), 
            .I2(n616), .I3(n17127), .O(n841_adj_2178[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_563_6_lut (.I0(GND_net), .I1(n835_adj_2172[3]), 
            .I2(n595), .I3(n17041), .O(n834[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_21 (.CI(n17295), .I0(Product1_mul_temp[21]), .I1(GND_net), 
            .CO(n17296));
    SB_CARRY Alpha_15__I_0_11_add_570_12 (.CI(n17127), .I0(n842_adj_2179[9]), 
            .I1(n616), .CO(n17128));
    SB_CARRY Beta_15__I_0_add_570_8 (.CI(n16940), .I0(n842[5]), .I1(n616), 
            .CO(n16941));
    SB_CARRY Beta_15__I_0_add_569_9 (.CI(n16954), .I0(n841[6]), .I1(n613), 
            .CO(n16955));
    SB_CARRY add_1232_10 (.CI(n16908), .I0(n840[14]), .I1(n767_adj_2041), 
            .CO(n16909));
    SB_CARRY Beta_15__I_0_add_572_6 (.CI(n16918), .I0(n844[3]), .I1(n622), 
            .CO(n16919));
    SB_LUT4 Beta_15__I_0_add_572_5_lut (.I0(GND_net), .I1(n844[2]), .I2(n622), 
            .I3(n16917), .O(n843[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_20_lut (.I0(GND_net), .I1(Product1_mul_temp[20]), .I2(GND_net), 
            .I3(n17294), .O(\dCurrent[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_6_lut (.I0(GND_net), .I1(n840[3]), .I2(n610), 
            .I3(n16966), .O(n839[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_20 (.CI(n17294), .I0(Product1_mul_temp[20]), .I1(GND_net), 
            .CO(n17295));
    SB_LUT4 Alpha_15__I_0_11_add_570_11_lut (.I0(GND_net), .I1(n842_adj_2179[8]), 
            .I2(n616), .I3(n17126), .O(n841_adj_2178[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_5 (.CI(n16980), .I0(n839[2]), .I1(n607), 
            .CO(n16981));
    SB_LUT4 Beta_15__I_0_add_567_4_lut (.I0(GND_net), .I1(n839[1]), .I2(n607), 
            .I3(n16979), .O(n838_adj_2170[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_19_lut (.I0(GND_net), .I1(Product1_mul_temp[19]), .I2(GND_net), 
            .I3(n17293), .O(\dCurrent[21] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_19 (.CI(n17293), .I0(Product1_mul_temp[19]), .I1(GND_net), 
            .CO(n17294));
    SB_CARRY Beta_15__I_0_add_561_5 (.CI(n17070), .I0(n833[2]), .I1(dCurrent[2]), 
            .CO(n17071));
    SB_LUT4 add_8094_18_lut (.I0(GND_net), .I1(Product1_mul_temp[18]), .I2(GND_net), 
            .I3(n17292), .O(\dCurrent[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_11 (.CI(n17126), .I0(n842_adj_2179[8]), 
            .I1(n616), .CO(n17127));
    SB_CARRY add_8094_18 (.CI(n17292), .I0(Product1_mul_temp[18]), .I1(GND_net), 
            .CO(n17293));
    SB_LUT4 Alpha_15__I_0_11_add_570_10_lut (.I0(GND_net), .I1(n842_adj_2179[7]), 
            .I2(n616), .I3(n17125), .O(n841_adj_2178[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_17_lut (.I0(GND_net), .I1(Product1_mul_temp[17]), .I2(GND_net), 
            .I3(n17291), .O(\dCurrent[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_17 (.CI(n17291), .I0(Product1_mul_temp[17]), .I1(GND_net), 
            .CO(n17292));
    SB_LUT4 add_8094_16_lut (.I0(GND_net), .I1(Product1_mul_temp[16]), .I2(GND_net), 
            .I3(n17290), .O(\dCurrent[18] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_10 (.CI(n17125), .I0(n842_adj_2179[7]), 
            .I1(n616), .CO(n17126));
    SB_LUT4 add_1232_9_lut (.I0(GND_net), .I1(n839[14]), .I2(n763_adj_2054), 
            .I3(n16907), .O(Product4_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_9 (.CI(n16907), .I0(n839[14]), .I1(n763_adj_2054), 
            .CO(n16908));
    SB_CARRY add_8094_16 (.CI(n17290), .I0(Product1_mul_temp[16]), .I1(GND_net), 
            .CO(n17291));
    SB_LUT4 Alpha_15__I_0_11_add_570_9_lut (.I0(GND_net), .I1(n842_adj_2179[6]), 
            .I2(n616), .I3(n17124), .O(n841_adj_2178[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_9 (.CI(n17124), .I0(n842_adj_2179[6]), 
            .I1(n616), .CO(n17125));
    SB_CARRY Beta_15__I_0_add_572_5 (.CI(n16917), .I0(n844[2]), .I1(n622), 
            .CO(n16918));
    SB_LUT4 Alpha_15__I_0_11_add_570_8_lut (.I0(GND_net), .I1(n842_adj_2179[5]), 
            .I2(n616), .I3(n17123), .O(n841_adj_2178[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_6 (.CI(n16927), .I0(n843[3]), .I1(n619), 
            .CO(n16928));
    SB_LUT4 Beta_15__I_0_add_570_7_lut (.I0(GND_net), .I1(n842[4]), .I2(n616), 
            .I3(n16939), .O(n841[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_5_lut (.I0(GND_net), .I1(n843[2]), .I2(n619), 
            .I3(n16926), .O(n842[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_7 (.CI(n16939), .I0(n842[4]), .I1(n616), 
            .CO(n16940));
    SB_LUT4 Beta_15__I_0_add_570_6_lut (.I0(GND_net), .I1(n842[3]), .I2(n616), 
            .I3(n16938), .O(n841[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_566_3_lut (.I0(GND_net), .I1(n838_adj_2170[0]), 
            .I2(n604), .I3(n16993), .O(n837_adj_2171[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_15_lut (.I0(GND_net), .I1(Product1_mul_temp[15]), .I2(GND_net), 
            .I3(n17289), .O(\dCurrent[17] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_3 (.CI(n16993), .I0(n838_adj_2170[0]), 
            .I1(n604), .CO(n16994));
    SB_CARRY add_8094_15 (.CI(n17289), .I0(Product1_mul_temp[15]), .I1(GND_net), 
            .CO(n17290));
    SB_CARRY Beta_15__I_0_add_566_16 (.CI(n17006), .I0(n838_adj_2170[13]), 
            .I1(n757), .CO(n759));
    SB_LUT4 Beta_15__I_0_add_569_8_lut (.I0(GND_net), .I1(n841[5]), .I2(n613), 
            .I3(n16953), .O(n840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_8 (.CI(n16953), .I0(n841[5]), .I1(n613), 
            .CO(n16954));
    SB_LUT4 add_8094_14_lut (.I0(GND_net), .I1(Product1_mul_temp[14]), .I2(GND_net), 
            .I3(n17288), .O(\dCurrent[16] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_8 (.CI(n17123), .I0(n842_adj_2179[5]), 
            .I1(n616), .CO(n17124));
    SB_LUT4 Alpha_15__I_0_11_add_570_7_lut (.I0(GND_net), .I1(n842_adj_2179[4]), 
            .I2(n616), .I3(n17122), .O(n841_adj_2178[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_15 (.CI(n17020), .I0(n837_adj_2171[12]), 
            .I1(n601), .CO(n17021));
    SB_LUT4 Beta_15__I_0_add_569_7_lut (.I0(GND_net), .I1(n841[4]), .I2(n613), 
            .I3(n16952), .O(n840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_6 (.CI(n16966), .I0(n840[3]), .I1(n610), 
            .CO(n16967));
    SB_CARRY Beta_15__I_0_add_567_4 (.CI(n16979), .I0(n839[1]), .I1(n607), 
            .CO(n16980));
    SB_LUT4 Beta_15__I_0_add_568_5_lut (.I0(GND_net), .I1(n840[2]), .I2(n610), 
            .I3(n16965), .O(n839[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_3_lut (.I0(GND_net), .I1(n839[0]), .I2(n607), 
            .I3(n16978), .O(n838_adj_2170[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_3 (.CI(n16978), .I0(n839[0]), .I1(n607), 
            .CO(n16979));
    SB_LUT4 Beta_15__I_0_add_565_14_lut (.I0(GND_net), .I1(n837_adj_2171[11]), 
            .I2(n601), .I3(n17019), .O(n836[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_14 (.CI(n17288), .I0(Product1_mul_temp[14]), .I1(GND_net), 
            .CO(n17289));
    SB_CARRY Alpha_15__I_0_11_add_570_7 (.CI(n17122), .I0(n842_adj_2179[4]), 
            .I1(n616), .CO(n17123));
    SB_LUT4 add_8094_13_lut (.I0(GND_net), .I1(Product1_mul_temp[13]), .I2(GND_net), 
            .I3(n17287), .O(\dCurrent[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_570_6_lut (.I0(GND_net), .I1(n842_adj_2179[3]), 
            .I2(n616), .I3(n17121), .O(n841_adj_2178[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_566_2_lut (.I0(GND_net), .I1(n607), .I2(n604), 
            .I3(GND_net), .O(n837_adj_2171[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_566_15_lut (.I0(GND_net), .I1(n838_adj_2170[12]), 
            .I2(n604), .I3(n17005), .O(n837_adj_2171[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_14 (.CI(n17019), .I0(n837_adj_2171[11]), 
            .I1(n601), .CO(n17020));
    SB_LUT4 Beta_15__I_0_add_565_13_lut (.I0(GND_net), .I1(n837_adj_2171[10]), 
            .I2(n601), .I3(n17018), .O(n836[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_13 (.CI(n17287), .I0(Product1_mul_temp[13]), .I1(GND_net), 
            .CO(n17288));
    SB_CARRY Beta_15__I_0_add_566_15 (.CI(n17005), .I0(n838_adj_2170[12]), 
            .I1(n604), .CO(n17006));
    SB_LUT4 add_8094_12_lut (.I0(GND_net), .I1(Product1_mul_temp[12]), .I2(GND_net), 
            .I3(n17286), .O(\dCurrent[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_6 (.CI(n17121), .I0(n842_adj_2179[3]), 
            .I1(n616), .CO(n17122));
    SB_CARRY Beta_15__I_0_add_563_6 (.CI(n17041), .I0(n835_adj_2172[3]), 
            .I1(n595), .CO(n17042));
    SB_LUT4 Beta_15__I_0_add_561_4_lut (.I0(GND_net), .I1(n833[1]), .I2(dCurrent[2]), 
            .I3(n17069), .O(Product4_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_570_5_lut (.I0(GND_net), .I1(n842_adj_2179[2]), 
            .I2(n616), .I3(n17120), .O(n841_adj_2178[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_5 (.CI(n17120), .I0(n842_adj_2179[2]), 
            .I1(n616), .CO(n17121));
    SB_CARRY add_8094_12 (.CI(n17286), .I0(Product1_mul_temp[12]), .I1(GND_net), 
            .CO(n17287));
    SB_LUT4 add_8094_11_lut (.I0(GND_net), .I1(Product1_mul_temp[11]), .I2(GND_net), 
            .I3(n17285), .O(\dCurrent[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_11 (.CI(n17285), .I0(Product1_mul_temp[11]), .I1(GND_net), 
            .CO(n17286));
    SB_LUT4 Alpha_15__I_0_11_add_570_4_lut (.I0(GND_net), .I1(n842_adj_2179[1]), 
            .I2(n616), .I3(n17119), .O(n841_adj_2178[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_10_lut (.I0(GND_net), .I1(Product1_mul_temp[10]), .I2(GND_net), 
            .I3(n17284), .O(\dCurrent[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_10 (.CI(n17284), .I0(Product1_mul_temp[10]), .I1(GND_net), 
            .CO(n17285));
    SB_LUT4 add_8094_9_lut (.I0(GND_net), .I1(Product1_mul_temp[9]), .I2(GND_net), 
            .I3(n17283), .O(\dCurrent[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_9 (.CI(n17283), .I0(Product1_mul_temp[9]), .I1(GND_net), 
            .CO(n17284));
    SB_LUT4 add_8094_8_lut (.I0(GND_net), .I1(Product1_mul_temp[8]), .I2(GND_net), 
            .I3(n17282), .O(\dCurrent[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_13 (.CI(n17018), .I0(n837_adj_2171[10]), 
            .I1(n601), .CO(n17019));
    SB_CARRY add_8094_8 (.CI(n17282), .I0(Product1_mul_temp[8]), .I1(GND_net), 
            .CO(n17283));
    SB_LUT4 add_8094_7_lut (.I0(GND_net), .I1(Product1_mul_temp[7]), .I2(GND_net), 
            .I3(n17281), .O(\dCurrent[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_7 (.CI(n17281), .I0(Product1_mul_temp[7]), .I1(GND_net), 
            .CO(n17282));
    SB_LUT4 add_8094_6_lut (.I0(GND_net), .I1(Product1_mul_temp[6]), .I2(GND_net), 
            .I3(n17280), .O(\dCurrent[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_563_5_lut (.I0(GND_net), .I1(n835_adj_2172[2]), 
            .I2(n595), .I3(n17040), .O(n834[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_6 (.CI(n17280), .I0(Product1_mul_temp[6]), .I1(GND_net), 
            .CO(n17281));
    SB_LUT4 add_8094_5_lut (.I0(GND_net), .I1(Product1_mul_temp[5]), .I2(GND_net), 
            .I3(n17279), .O(\dCurrent[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_5 (.CI(n17279), .I0(Product1_mul_temp[5]), .I1(GND_net), 
            .CO(n17280));
    SB_CARRY Beta_15__I_0_add_566_2 (.CI(GND_net), .I0(n607), .I1(n604), 
            .CO(n16993));
    SB_LUT4 add_8094_4_lut (.I0(GND_net), .I1(Product1_mul_temp[4]), .I2(GND_net), 
            .I3(n17278), .O(\dCurrent[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_4 (.CI(n17069), .I0(n833[1]), .I1(dCurrent[2]), 
            .CO(n17070));
    SB_LUT4 Beta_15__I_0_add_567_16_lut (.I0(GND_net), .I1(n839[13]), .I2(n761), 
            .I3(n16991), .O(n838_adj_2170[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_4 (.CI(n17278), .I0(Product1_mul_temp[4]), .I1(GND_net), 
            .CO(n17279));
    SB_CARRY Alpha_15__I_0_11_add_570_4 (.CI(n17119), .I0(n842_adj_2179[1]), 
            .I1(n616), .CO(n17120));
    SB_LUT4 add_8094_3_lut (.I0(GND_net), .I1(Product1_mul_temp[3]), .I2(GND_net), 
            .I3(n17277), .O(\dCurrent[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_3 (.CI(n17277), .I0(Product1_mul_temp[3]), .I1(GND_net), 
            .CO(n17278));
    SB_LUT4 Beta_15__I_0_add_566_14_lut (.I0(GND_net), .I1(n838_adj_2170[11]), 
            .I2(n604), .I3(n17004), .O(n837_adj_2171[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_570_3_lut (.I0(GND_net), .I1(n842_adj_2179[0]), 
            .I2(n616), .I3(n17118), .O(n841_adj_2178[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_8094_2_lut (.I0(GND_net), .I1(Product1_mul_temp[2]), .I2(\Product_mul_temp[26] ), 
            .I3(GND_net), .O(\dCurrent[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_8094_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_8094_2 (.CI(GND_net), .I0(Product1_mul_temp[2]), .I1(\Product_mul_temp[26] ), 
            .CO(n17277));
    SB_LUT4 Beta_15__I_0_add_565_12_lut (.I0(GND_net), .I1(n837_adj_2171[9]), 
            .I2(n601), .I3(n17017), .O(n836[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_5 (.CI(n17040), .I0(n835_adj_2172[2]), 
            .I1(n595), .CO(n17041));
    SB_LUT4 Beta_15__I_0_add_563_4_lut (.I0(GND_net), .I1(n835_adj_2172[1]), 
            .I2(n595), .I3(n17039), .O(n834[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_3 (.CI(n17118), .I0(n842_adj_2179[0]), 
            .I1(n616), .CO(n17119));
    SB_CARRY Beta_15__I_0_add_563_4 (.CI(n17039), .I0(n835_adj_2172[1]), 
            .I1(n595), .CO(n17040));
    SB_LUT4 Alpha_15__I_0_11_add_570_2_lut (.I0(GND_net), .I1(n619), .I2(n616), 
            .I3(GND_net), .O(n841_adj_2178[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_561_3_lut (.I0(GND_net), .I1(n833[0]), .I2(dCurrent[2]), 
            .I3(n17068), .O(Product4_mul_temp[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_570_2 (.CI(GND_net), .I0(n619), .I1(n616), 
            .CO(n17118));
    SB_CARRY Beta_15__I_0_add_561_3 (.CI(n17068), .I0(n833[0]), .I1(dCurrent[2]), 
            .CO(n17069));
    SB_LUT4 Alpha_15__I_0_11_add_571_12_lut (.I0(GND_net), .I1(n843_adj_2180[7]), 
            .I2(n777), .I3(n17116), .O(n842_adj_2179[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_571_12 (.CI(n17116), .I0(n843_adj_2180[7]), 
            .I1(n777), .CO(n779_adj_2070));
    SB_LUT4 Beta_15__I_0_add_561_2_lut (.I0(GND_net), .I1(n592), .I2(dCurrent[2]), 
            .I3(GND_net), .O(\qCurrent[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_561_16_lut (.I0(GND_net), .I1(n833_adj_2175[13]), 
            .I2(n737), .I3(n17264), .O(n832[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_16 (.CI(n17264), .I0(n833_adj_2175[13]), 
            .I1(n737), .CO(n739));
    SB_LUT4 Alpha_15__I_0_11_add_561_15_lut (.I0(GND_net), .I1(n833_adj_2175[12]), 
            .I2(dCurrent[2]), .I3(n17263), .O(Product1_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_571_11_lut (.I0(GND_net), .I1(n843_adj_2180[7]), 
            .I2(n619), .I3(n17115), .O(n842_adj_2179[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_15 (.CI(n17263), .I0(n833_adj_2175[12]), 
            .I1(dCurrent[2]), .CO(n17264));
    SB_LUT4 Alpha_15__I_0_11_add_561_14_lut (.I0(GND_net), .I1(n833_adj_2175[11]), 
            .I2(dCurrent[2]), .I3(n17262), .O(Product1_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_14 (.CI(n17262), .I0(n833_adj_2175[11]), 
            .I1(dCurrent[2]), .CO(n17263));
    SB_LUT4 Alpha_15__I_0_11_add_561_13_lut (.I0(GND_net), .I1(n833_adj_2175[10]), 
            .I2(dCurrent[2]), .I3(n17261), .O(Product1_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1232_8_lut (.I0(GND_net), .I1(n838_adj_2170[14]), .I2(n759), 
            .I3(n16906), .O(Product4_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_8 (.CI(n16906), .I0(n838_adj_2170[14]), .I1(n759), 
            .CO(n16907));
    SB_CARRY Alpha_15__I_0_11_add_561_13 (.CI(n17261), .I0(n833_adj_2175[10]), 
            .I1(dCurrent[2]), .CO(n17262));
    SB_CARRY Alpha_15__I_0_11_add_571_11 (.CI(n17115), .I0(n843_adj_2180[7]), 
            .I1(n619), .CO(n17116));
    SB_LUT4 Beta_15__I_0_add_572_4_lut (.I0(GND_net), .I1(n844[1]), .I2(n622), 
            .I3(n16916), .O(n843[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_5 (.CI(n16926), .I0(n843[2]), .I1(n619), 
            .CO(n16927));
    SB_CARRY Beta_15__I_0_add_570_6 (.CI(n16938), .I0(n842[3]), .I1(n616), 
            .CO(n16939));
    SB_LUT4 Beta_15__I_0_add_570_5_lut (.I0(GND_net), .I1(n842[2]), .I2(n616), 
            .I3(n16937), .O(n841[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_561_12_lut (.I0(GND_net), .I1(n833_adj_2175[9]), 
            .I2(dCurrent[2]), .I3(n17260), .O(Product1_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_571_10_lut (.I0(GND_net), .I1(n843_adj_2180[7]), 
            .I2(n619), .I3(n17114), .O(n842_adj_2179[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_7 (.CI(n16952), .I0(n841[4]), .I1(n613), 
            .CO(n16953));
    SB_CARRY Beta_15__I_0_add_568_5 (.CI(n16965), .I0(n840[2]), .I1(n610), 
            .CO(n16966));
    SB_LUT4 Beta_15__I_0_add_567_2_lut (.I0(GND_net), .I1(n610), .I2(n607), 
            .I3(GND_net), .O(n838_adj_2170[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_2 (.CI(GND_net), .I0(n610), .I1(n607), 
            .CO(n16978));
    SB_CARRY Alpha_15__I_0_11_add_561_12 (.CI(n17260), .I0(n833_adj_2175[9]), 
            .I1(dCurrent[2]), .CO(n17261));
    SB_CARRY Alpha_15__I_0_11_add_571_10 (.CI(n17114), .I0(n843_adj_2180[7]), 
            .I1(n619), .CO(n17115));
    SB_CARRY Beta_15__I_0_add_567_16 (.CI(n16991), .I0(n839[13]), .I1(n761), 
            .CO(n763_adj_2054));
    SB_CARRY Beta_15__I_0_add_566_14 (.CI(n17004), .I0(n838_adj_2170[11]), 
            .I1(n604), .CO(n17005));
    SB_LUT4 Beta_15__I_0_add_566_13_lut (.I0(GND_net), .I1(n838_adj_2170[10]), 
            .I2(n604), .I3(n17003), .O(n837_adj_2171[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_2 (.CI(GND_net), .I0(n592), .I1(dCurrent[2]), 
            .CO(n17068));
    SB_LUT4 Alpha_15__I_0_11_add_571_9_lut (.I0(GND_net), .I1(n843_adj_2180[6]), 
            .I2(n619), .I3(n17113), .O(n842_adj_2179[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_571_9 (.CI(n17113), .I0(n843_adj_2180[6]), 
            .I1(n619), .CO(n17114));
    SB_LUT4 Alpha_15__I_0_11_add_561_11_lut (.I0(GND_net), .I1(n833_adj_2175[8]), 
            .I2(dCurrent[2]), .I3(n17259), .O(Product1_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_11 (.CI(n17259), .I0(n833_adj_2175[8]), 
            .I1(dCurrent[2]), .CO(n17260));
    SB_LUT4 Alpha_15__I_0_11_add_571_8_lut (.I0(GND_net), .I1(n843_adj_2180[5]), 
            .I2(n619), .I3(n17112), .O(n842_adj_2179[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_571_8 (.CI(n17112), .I0(n843_adj_2180[5]), 
            .I1(n619), .CO(n17113));
    SB_LUT4 Alpha_15__I_0_11_add_561_10_lut (.I0(GND_net), .I1(n833_adj_2175[7]), 
            .I2(dCurrent[2]), .I3(n17258), .O(Product1_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_10 (.CI(n17258), .I0(n833_adj_2175[7]), 
            .I1(dCurrent[2]), .CO(n17259));
    SB_LUT4 Alpha_15__I_0_11_add_561_9_lut (.I0(GND_net), .I1(n833_adj_2175[6]), 
            .I2(dCurrent[2]), .I3(n17257), .O(Product1_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_9 (.CI(n17257), .I0(n833_adj_2175[6]), 
            .I1(dCurrent[2]), .CO(n17258));
    SB_LUT4 Alpha_15__I_0_11_add_561_8_lut (.I0(GND_net), .I1(n833_adj_2175[5]), 
            .I2(dCurrent[2]), .I3(n17256), .O(Product1_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_8 (.CI(n17256), .I0(n833_adj_2175[5]), 
            .I1(dCurrent[2]), .CO(n17257));
    SB_LUT4 Alpha_15__I_0_11_add_561_7_lut (.I0(GND_net), .I1(n833_adj_2175[4]), 
            .I2(dCurrent[2]), .I3(n17255), .O(Product1_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_7 (.CI(n17255), .I0(n833_adj_2175[4]), 
            .I1(dCurrent[2]), .CO(n17256));
    SB_LUT4 Alpha_15__I_0_11_add_561_6_lut (.I0(GND_net), .I1(n833_adj_2175[3]), 
            .I2(dCurrent[2]), .I3(n17254), .O(Product1_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_12 (.CI(n17017), .I0(n837_adj_2171[9]), 
            .I1(n601), .CO(n17018));
    SB_LUT4 Beta_15__I_0_add_563_3_lut (.I0(GND_net), .I1(n835_adj_2172[0]), 
            .I2(n595), .I3(n17038), .O(n834[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_16_lut (.I0(GND_net), .I1(n834[13]), .I2(n741), 
            .I3(n17066), .O(n833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_6 (.CI(n17254), .I0(n833_adj_2175[3]), 
            .I1(dCurrent[2]), .CO(n17255));
    SB_LUT4 Alpha_15__I_0_11_add_571_7_lut (.I0(GND_net), .I1(n843_adj_2180[4]), 
            .I2(n619), .I3(n17111), .O(n842_adj_2179[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1232_7_lut (.I0(GND_net), .I1(n837_adj_2171[14]), .I2(n755), 
            .I3(n16905), .O(Product4_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_4 (.CI(n16916), .I0(n844[1]), .I1(n622), 
            .CO(n16917));
    SB_LUT4 Beta_15__I_0_add_572_3_lut (.I0(GND_net), .I1(n844[0]), .I2(n622), 
            .I3(n16915), .O(n843[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_561_5_lut (.I0(GND_net), .I1(n833_adj_2175[2]), 
            .I2(dCurrent[2]), .I3(n17253), .O(Product1_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_571_7 (.CI(n17111), .I0(n843_adj_2180[4]), 
            .I1(n619), .CO(n17112));
    SB_LUT4 Beta_15__I_0_add_571_4_lut (.I0(GND_net), .I1(n843[1]), .I2(n619), 
            .I3(n16925), .O(n842[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_5 (.CI(n16937), .I0(n842[2]), .I1(n616), 
            .CO(n16938));
    SB_LUT4 Beta_15__I_0_add_569_6_lut (.I0(GND_net), .I1(n841[3]), .I2(n613), 
            .I3(n16951), .O(n840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_6 (.CI(n16951), .I0(n841[3]), .I1(n613), 
            .CO(n16952));
    SB_CARRY Alpha_15__I_0_11_add_561_5 (.CI(n17253), .I0(n833_adj_2175[2]), 
            .I1(dCurrent[2]), .CO(n17254));
    SB_LUT4 Alpha_15__I_0_11_add_571_6_lut (.I0(GND_net), .I1(n843_adj_2180[3]), 
            .I2(n619), .I3(n17110), .O(n842_adj_2179[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_4_lut (.I0(GND_net), .I1(n840[1]), .I2(n610), 
            .I3(n16964), .O(n839[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_16_lut (.I0(GND_net), .I1(n840[13]), .I2(n765), 
            .I3(n16976), .O(n839[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_15_lut (.I0(GND_net), .I1(n839[12]), .I2(n607), 
            .I3(n16990), .O(n838_adj_2170[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_15 (.CI(n16990), .I0(n839[12]), .I1(n607), 
            .CO(n16991));
    SB_LUT4 Alpha_15__I_0_11_add_561_4_lut (.I0(GND_net), .I1(n833_adj_2175[1]), 
            .I2(dCurrent[2]), .I3(n17252), .O(Product1_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_571_6 (.CI(n17110), .I0(n843_adj_2180[3]), 
            .I1(n619), .CO(n17111));
    SB_CARRY Beta_15__I_0_add_566_13 (.CI(n17003), .I0(n838_adj_2170[10]), 
            .I1(n604), .CO(n17004));
    SB_LUT4 Beta_15__I_0_add_565_11_lut (.I0(GND_net), .I1(n837_adj_2171[8]), 
            .I2(n601), .I3(n17016), .O(n836[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_3 (.CI(n17038), .I0(n835_adj_2172[0]), 
            .I1(n595), .CO(n17039));
    SB_LUT4 Beta_15__I_0_add_563_2_lut (.I0(GND_net), .I1(n598), .I2(n595), 
            .I3(GND_net), .O(n834[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_571_5_lut (.I0(GND_net), .I1(n843_adj_2180[2]), 
            .I2(n619), .I3(n17109), .O(n842_adj_2179[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_4 (.CI(n17252), .I0(n833_adj_2175[1]), 
            .I1(dCurrent[2]), .CO(n17253));
    SB_LUT4 Alpha_15__I_0_11_add_561_3_lut (.I0(GND_net), .I1(n833_adj_2175[0]), 
            .I2(dCurrent[2]), .I3(n17251), .O(Product1_mul_temp[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_571_5 (.CI(n17109), .I0(n843_adj_2180[2]), 
            .I1(n619), .CO(n17110));
    SB_LUT4 Beta_15__I_0_i519_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n765));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i519_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY Alpha_15__I_0_11_add_561_3 (.CI(n17251), .I0(n833_adj_2175[0]), 
            .I1(dCurrent[2]), .CO(n17252));
    SB_LUT4 Alpha_15__I_0_11_add_561_2_lut (.I0(GND_net), .I1(n592), .I2(dCurrent[2]), 
            .I3(GND_net), .O(\dCurrent[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_561_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_561_2 (.CI(GND_net), .I0(n592), .I1(dCurrent[2]), 
            .CO(n17251));
    SB_CARRY Beta_15__I_0_add_562_16 (.CI(n17066), .I0(n834[13]), .I1(n741), 
            .CO(n743_adj_2096));
    SB_LUT4 Alpha_15__I_0_11_add_562_16_lut (.I0(GND_net), .I1(n834_adj_2173[13]), 
            .I2(n741), .I3(n17249), .O(n833_adj_2175[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_16 (.CI(n17249), .I0(n834_adj_2173[13]), 
            .I1(n741), .CO(n743));
    SB_LUT4 Alpha_15__I_0_11_add_562_15_lut (.I0(GND_net), .I1(n834_adj_2173[12]), 
            .I2(n592), .I3(n17248), .O(n833_adj_2175[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_15 (.CI(n17248), .I0(n834_adj_2173[12]), 
            .I1(n592), .CO(n17249));
    SB_LUT4 Alpha_15__I_0_11_add_562_14_lut (.I0(GND_net), .I1(n834_adj_2173[11]), 
            .I2(n592), .I3(n17247), .O(n833_adj_2175[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_14 (.CI(n17247), .I0(n834_adj_2173[11]), 
            .I1(n592), .CO(n17248));
    SB_LUT4 Alpha_15__I_0_11_add_562_13_lut (.I0(GND_net), .I1(n834_adj_2173[10]), 
            .I2(n592), .I3(n17246), .O(n833_adj_2175[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_15_lut (.I0(GND_net), .I1(n834[12]), .I2(n592), 
            .I3(n17065), .O(n833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_571_4_lut (.I0(GND_net), .I1(n843_adj_2180[1]), 
            .I2(n619), .I3(n17108), .O(n842_adj_2179[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_13 (.CI(n17246), .I0(n834_adj_2173[10]), 
            .I1(n592), .CO(n17247));
    SB_LUT4 Alpha_15__I_0_11_i20_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n616));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Alpha_15__I_0_11_add_562_12_lut (.I0(GND_net), .I1(n834_adj_2173[9]), 
            .I2(n592), .I3(n17245), .O(n833_adj_2175[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_12 (.CI(n17245), .I0(n834_adj_2173[9]), 
            .I1(n592), .CO(n17246));
    SB_CARRY Alpha_15__I_0_11_add_571_4 (.CI(n17108), .I0(n843_adj_2180[1]), 
            .I1(n619), .CO(n17109));
    SB_LUT4 Beta_15__I_0_i507_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i507_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Alpha_15__I_0_11_add_562_11_lut (.I0(GND_net), .I1(n834_adj_2173[8]), 
            .I2(n592), .I3(n17244), .O(n833_adj_2175[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_571_3_lut (.I0(GND_net), .I1(n843_adj_2180[0]), 
            .I2(n619), .I3(n17107), .O(n842_adj_2179[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_i26_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n625));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_1232_7 (.CI(n16905), .I0(n837_adj_2171[14]), .I1(n755), 
            .CO(n16906));
    SB_LUT4 add_1232_6_lut (.I0(GND_net), .I1(n836[14]), .I2(n751), .I3(n16904), 
            .O(Product4_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_11 (.CI(n17244), .I0(n834_adj_2173[8]), 
            .I1(n592), .CO(n17245));
    SB_CARRY Alpha_15__I_0_11_add_571_3 (.CI(n17107), .I0(n843_adj_2180[0]), 
            .I1(n619), .CO(n17108));
    SB_CARRY Beta_15__I_0_add_572_3 (.CI(n16915), .I0(n844[0]), .I1(n622), 
            .CO(n16916));
    SB_CARRY Beta_15__I_0_add_571_4 (.CI(n16925), .I0(n843[1]), .I1(n619), 
            .CO(n16926));
    SB_LUT4 Beta_15__I_0_add_570_4_lut (.I0(GND_net), .I1(n842[1]), .I2(n616), 
            .I3(n16936), .O(n841[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_4 (.CI(n16936), .I0(n842[1]), .I1(n616), 
            .CO(n16937));
    SB_LUT4 Alpha_15__I_0_11_add_562_10_lut (.I0(GND_net), .I1(n834_adj_2173[7]), 
            .I2(n592), .I3(n17243), .O(n833_adj_2175[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_571_2_lut (.I0(GND_net), .I1(n622), .I2(n619), 
            .I3(GND_net), .O(n842_adj_2179[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_5_lut (.I0(GND_net), .I1(n841[2]), .I2(n613), 
            .I3(n16950), .O(n840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_4 (.CI(n16964), .I0(n840[1]), .I1(n610), 
            .CO(n16965));
    SB_CARRY Beta_15__I_0_add_568_16 (.CI(n16976), .I0(n840[13]), .I1(n765), 
            .CO(n767_adj_2041));
    SB_LUT4 Beta_15__I_0_add_568_15_lut (.I0(GND_net), .I1(n840[12]), .I2(n610), 
            .I3(n16975), .O(n839[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_i531_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n781));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i531_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY Alpha_15__I_0_11_add_562_10 (.CI(n17243), .I0(n834_adj_2173[7]), 
            .I1(n592), .CO(n17244));
    SB_CARRY Alpha_15__I_0_11_add_571_2 (.CI(GND_net), .I0(n622), .I1(n619), 
            .CO(n17107));
    SB_LUT4 Beta_15__I_0_add_567_14_lut (.I0(GND_net), .I1(n839[11]), .I2(n607), 
            .I3(n16989), .O(n838_adj_2170[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_566_12_lut (.I0(GND_net), .I1(n838_adj_2170[9]), 
            .I2(n604), .I3(n17002), .O(n837_adj_2171[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_11 (.CI(n17016), .I0(n837_adj_2171[8]), 
            .I1(n601), .CO(n17017));
    SB_LUT4 Beta_15__I_0_add_565_10_lut (.I0(GND_net), .I1(n837_adj_2171[7]), 
            .I2(n601), .I3(n17015), .O(n836[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_562_9_lut (.I0(GND_net), .I1(n834_adj_2173[6]), 
            .I2(n592), .I3(n17242), .O(n833_adj_2175[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_15 (.CI(n17065), .I0(n834[12]), .I1(n592), 
            .CO(n17066));
    SB_LUT4 Alpha_15__I_0_11_add_572_10_lut (.I0(GND_net), .I1(n844_adj_2181[5]), 
            .I2(n781), .I3(n17105), .O(n843_adj_2180[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_572_10 (.CI(n17105), .I0(n844_adj_2181[5]), 
            .I1(n781), .CO(n783));
    SB_CARRY Alpha_15__I_0_11_add_562_9 (.CI(n17242), .I0(n834_adj_2173[6]), 
            .I1(n592), .CO(n17243));
    SB_LUT4 Alpha_15__I_0_11_add_562_8_lut (.I0(GND_net), .I1(n834_adj_2173[5]), 
            .I2(n592), .I3(n17241), .O(n833_adj_2175[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_572_9_lut (.I0(GND_net), .I1(n844_adj_2181[5]), 
            .I2(n622), .I3(n17104), .O(n843_adj_2180[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_8 (.CI(n17241), .I0(n834_adj_2173[5]), 
            .I1(n592), .CO(n17242));
    SB_LUT4 Alpha_15__I_0_11_add_562_7_lut (.I0(GND_net), .I1(n834_adj_2173[4]), 
            .I2(n592), .I3(n17240), .O(n833_adj_2175[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_7 (.CI(n17240), .I0(n834_adj_2173[4]), 
            .I1(n592), .CO(n17241));
    SB_LUT4 Alpha_15__I_0_11_add_562_6_lut (.I0(GND_net), .I1(n834_adj_2173[3]), 
            .I2(n592), .I3(n17239), .O(n833_adj_2175[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_6 (.CI(n17239), .I0(n834_adj_2173[3]), 
            .I1(n592), .CO(n17240));
    SB_LUT4 Alpha_15__I_0_11_add_562_5_lut (.I0(GND_net), .I1(n834_adj_2173[2]), 
            .I2(n592), .I3(n17238), .O(n833_adj_2175[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_5 (.CI(n17238), .I0(n834_adj_2173[2]), 
            .I1(n592), .CO(n17239));
    SB_LUT4 Alpha_15__I_0_11_add_562_4_lut (.I0(GND_net), .I1(n834_adj_2173[1]), 
            .I2(n592), .I3(n17237), .O(n833_adj_2175[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_4 (.CI(n17237), .I0(n834_adj_2173[1]), 
            .I1(n592), .CO(n17238));
    SB_CARRY Beta_15__I_0_add_563_2 (.CI(GND_net), .I0(n598), .I1(n595), 
            .CO(n17038));
    SB_LUT4 Beta_15__I_0_add_562_14_lut (.I0(GND_net), .I1(n834[11]), .I2(n592), 
            .I3(n17064), .O(n833[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_14 (.CI(n17064), .I0(n834[11]), .I1(n592), 
            .CO(n17065));
    SB_LUT4 Alpha_15__I_0_11_add_562_3_lut (.I0(GND_net), .I1(n834_adj_2173[0]), 
            .I2(n592), .I3(n17236), .O(n833_adj_2175[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_3 (.CI(n17236), .I0(n834_adj_2173[0]), 
            .I1(n592), .CO(n17237));
    SB_LUT4 Alpha_15__I_0_11_i24_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n622));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Beta_15__I_0_i504_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n745));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i504_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Beta_15__I_0_i501_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n741));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i501_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY Alpha_15__I_0_11_add_572_9 (.CI(n17104), .I0(n844_adj_2181[5]), 
            .I1(n622), .CO(n17105));
    SB_LUT4 Alpha_15__I_0_11_add_562_2_lut (.I0(GND_net), .I1(n595), .I2(n592), 
            .I3(GND_net), .O(n833_adj_2175[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_572_8_lut (.I0(GND_net), .I1(n844_adj_2181[5]), 
            .I2(n622), .I3(n17103), .O(n843_adj_2180[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_6 (.CI(n16904), .I0(n836[14]), .I1(n751), .CO(n16905));
    SB_LUT4 add_1232_5_lut (.I0(GND_net), .I1(n835_adj_2172[14]), .I2(n747_adj_2012), 
            .I3(n16903), .O(Product4_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_562_2 (.CI(GND_net), .I0(n595), .I1(n592), 
            .CO(n17236));
    SB_CARRY Alpha_15__I_0_11_add_572_8 (.CI(n17103), .I0(n844_adj_2181[5]), 
            .I1(n622), .CO(n17104));
    SB_LUT4 Beta_15__I_0_add_572_2_lut (.I0(GND_net), .I1(n625), .I2(n622), 
            .I3(GND_net), .O(n843[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_3_lut (.I0(GND_net), .I1(n843[0]), .I2(n619), 
            .I3(n16924), .O(n842[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_3_lut (.I0(GND_net), .I1(n842[0]), .I2(n616), 
            .I3(n16935), .O(n841[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_3 (.CI(n16935), .I0(n842[0]), .I1(n616), 
            .CO(n16936));
    SB_LUT4 Alpha_15__I_0_11_add_563_16_lut (.I0(GND_net), .I1(n835[13]), 
            .I2(n745), .I3(n17234), .O(n834_adj_2173[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_572_7_lut (.I0(GND_net), .I1(n844_adj_2181[4]), 
            .I2(n622), .I3(n17102), .O(n843_adj_2180[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_5 (.CI(n16950), .I0(n841[2]), .I1(n613), 
            .CO(n16951));
    SB_LUT4 Beta_15__I_0_add_568_3_lut (.I0(GND_net), .I1(n840[0]), .I2(n610), 
            .I3(n16963), .O(n839[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_15 (.CI(n16975), .I0(n840[12]), .I1(n610), 
            .CO(n16976));
    SB_LUT4 Beta_15__I_0_add_568_14_lut (.I0(GND_net), .I1(n840[11]), .I2(n610), 
            .I3(n16974), .O(n839[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_16 (.CI(n17234), .I0(n835[13]), .I1(n745), 
            .CO(n747));
    SB_CARRY Alpha_15__I_0_11_add_572_7 (.CI(n17102), .I0(n844_adj_2181[4]), 
            .I1(n622), .CO(n17103));
    SB_CARRY Beta_15__I_0_add_567_14 (.CI(n16989), .I0(n839[11]), .I1(n607), 
            .CO(n16990));
    SB_CARRY Beta_15__I_0_add_566_12 (.CI(n17002), .I0(n838_adj_2170[9]), 
            .I1(n604), .CO(n17003));
    SB_CARRY Beta_15__I_0_add_565_10 (.CI(n17015), .I0(n837_adj_2171[7]), 
            .I1(n601), .CO(n17016));
    SB_LUT4 Beta_15__I_0_add_565_9_lut (.I0(GND_net), .I1(n837_adj_2171[6]), 
            .I2(n601), .I3(n17014), .O(n836[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_563_15_lut (.I0(GND_net), .I1(n835[12]), 
            .I2(n595), .I3(n17233), .O(n834_adj_2173[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_572_6_lut (.I0(GND_net), .I1(n844_adj_2181[3]), 
            .I2(n622), .I3(n17101), .O(n843_adj_2180[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_16_lut (.I0(GND_net), .I1(n836[13]), .I2(n749), 
            .I3(n17036), .O(n835_adj_2172[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_13_lut (.I0(GND_net), .I1(n834[10]), .I2(n592), 
            .I3(n17063), .O(n833[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_572_6 (.CI(n17101), .I0(n844_adj_2181[3]), 
            .I1(n622), .CO(n17102));
    SB_LUT4 Alpha_15__I_0_11_add_572_5_lut (.I0(GND_net), .I1(n844_adj_2181[2]), 
            .I2(n622), .I3(n17100), .O(n843_adj_2180[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_i6_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n595));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Alpha_15__I_0_11_add_572_5 (.CI(n17100), .I0(n844_adj_2181[2]), 
            .I1(n622), .CO(n17101));
    SB_LUT4 Alpha_15__I_0_11_i2_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(dCurrent[2]));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Alpha_15__I_0_11_add_563_15 (.CI(n17233), .I0(n835[12]), .I1(n595), 
            .CO(n17234));
    SB_LUT4 Alpha_15__I_0_11_add_572_4_lut (.I0(GND_net), .I1(n844_adj_2181[1]), 
            .I2(n622), .I3(n17099), .O(n843_adj_2180[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_572_4 (.CI(n17099), .I0(n844_adj_2181[1]), 
            .I1(n622), .CO(n17100));
    SB_LUT4 Alpha_15__I_0_11_add_563_14_lut (.I0(GND_net), .I1(n835[11]), 
            .I2(n595), .I3(n17232), .O(n834_adj_2173[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_14 (.CI(n17232), .I0(n835[11]), .I1(n595), 
            .CO(n17233));
    SB_LUT4 Alpha_15__I_0_11_add_563_13_lut (.I0(GND_net), .I1(n835[10]), 
            .I2(n595), .I3(n17231), .O(n834_adj_2173[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_13 (.CI(n17231), .I0(n835[10]), .I1(n595), 
            .CO(n17232));
    SB_LUT4 Alpha_15__I_0_11_add_563_12_lut (.I0(GND_net), .I1(n835[9]), 
            .I2(n595), .I3(n17230), .O(n834_adj_2173[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_16 (.CI(n17036), .I0(n836[13]), .I1(n749), 
            .CO(n751));
    SB_CARRY Alpha_15__I_0_11_add_563_12 (.CI(n17230), .I0(n835[9]), .I1(n595), 
            .CO(n17231));
    SB_LUT4 Alpha_15__I_0_11_add_563_11_lut (.I0(GND_net), .I1(n835[8]), 
            .I2(n595), .I3(n17229), .O(n834_adj_2173[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_11 (.CI(n17229), .I0(n835[8]), .I1(n595), 
            .CO(n17230));
    SB_LUT4 Alpha_15__I_0_11_add_563_10_lut (.I0(GND_net), .I1(n835[7]), 
            .I2(n595), .I3(n17228), .O(n834_adj_2173[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_10 (.CI(n17228), .I0(n835[7]), .I1(n595), 
            .CO(n17229));
    SB_LUT4 Alpha_15__I_0_11_add_563_9_lut (.I0(GND_net), .I1(n835[6]), 
            .I2(n595), .I3(n17227), .O(n834_adj_2173[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_9 (.CI(n17227), .I0(n835[6]), .I1(n595), 
            .CO(n17228));
    SB_LUT4 Alpha_15__I_0_11_add_563_8_lut (.I0(GND_net), .I1(n835[5]), 
            .I2(n595), .I3(n17226), .O(n834_adj_2173[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_8 (.CI(n17226), .I0(n835[5]), .I1(n595), 
            .CO(n17227));
    SB_LUT4 Alpha_15__I_0_11_add_563_7_lut (.I0(GND_net), .I1(n835[4]), 
            .I2(n595), .I3(n17225), .O(n834_adj_2173[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_7 (.CI(n17225), .I0(n835[4]), .I1(n595), 
            .CO(n17226));
    SB_LUT4 Alpha_15__I_0_11_add_563_6_lut (.I0(GND_net), .I1(n835[3]), 
            .I2(n595), .I3(n17224), .O(n834_adj_2173[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_6 (.CI(n17224), .I0(n835[3]), .I1(n595), 
            .CO(n17225));
    SB_LUT4 Alpha_15__I_0_11_add_563_5_lut (.I0(GND_net), .I1(n835[2]), 
            .I2(n595), .I3(n17223), .O(n834_adj_2173[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_5 (.CI(n17223), .I0(n835[2]), .I1(n595), 
            .CO(n17224));
    SB_LUT4 Alpha_15__I_0_11_add_572_3_lut (.I0(GND_net), .I1(n844_adj_2181[0]), 
            .I2(n622), .I3(n17098), .O(n843_adj_2180[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_563_4_lut (.I0(GND_net), .I1(n835[1]), 
            .I2(n595), .I3(n17222), .O(n834_adj_2173[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_572_3 (.CI(n17098), .I0(n844_adj_2181[0]), 
            .I1(n622), .CO(n17099));
    SB_CARRY Alpha_15__I_0_11_add_563_4 (.CI(n17222), .I0(n835[1]), .I1(n595), 
            .CO(n17223));
    SB_LUT4 Beta_15__I_0_add_573_8_lut (.I0(GND_net), .I1(n845[3]), .I2(n785), 
            .I3(n18165), .O(n844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_8 (.CI(n18165), .I0(n845[3]), .I1(n785), 
            .CO(n787));
    SB_LUT4 Beta_15__I_0_add_573_7_lut (.I0(GND_net), .I1(n845[3]), .I2(n625), 
            .I3(n18164), .O(n844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_7 (.CI(n18164), .I0(n845[3]), .I1(n625), 
            .CO(n18165));
    SB_LUT4 Beta_15__I_0_add_573_6_lut (.I0(GND_net), .I1(n845[3]), .I2(n625), 
            .I3(n18163), .O(n844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_6 (.CI(n18163), .I0(n845[3]), .I1(n625), 
            .CO(n18164));
    SB_LUT4 Beta_15__I_0_add_573_5_lut (.I0(GND_net), .I1(n845[2]), .I2(n625), 
            .I3(n18162), .O(n844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_5 (.CI(n18162), .I0(n845[2]), .I1(n625), 
            .CO(n18163));
    SB_LUT4 Beta_15__I_0_add_573_4_lut (.I0(GND_net), .I1(n139), .I2(n625), 
            .I3(n18161), .O(n844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_4 (.CI(n18161), .I0(n139), .I1(n625), 
            .CO(n18162));
    SB_LUT4 Beta_15__I_0_add_573_3_lut (.I0(GND_net), .I1(n845[0]), .I2(n625), 
            .I3(n18160), .O(n844[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_3 (.CI(n18160), .I0(n845[0]), .I1(n625), 
            .CO(n18161));
    SB_LUT4 Beta_15__I_0_add_573_2_lut (.I0(GND_net), .I1(n628), .I2(n625), 
            .I3(GND_net), .O(n844[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_2 (.CI(GND_net), .I0(n628), .I1(n625), 
            .CO(n18160));
    SB_LUT4 Alpha_15__I_0_11_add_563_3_lut (.I0(GND_net), .I1(n835[0]), 
            .I2(n595), .I3(n17221), .O(n834_adj_2173[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_572_2_lut (.I0(GND_net), .I1(n625), .I2(n622), 
            .I3(GND_net), .O(n843_adj_2180[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_3 (.CI(n17221), .I0(n835[0]), .I1(n595), 
            .CO(n17222));
    SB_LUT4 Alpha_15__I_0_11_add_563_2_lut (.I0(GND_net), .I1(n598), .I2(n595), 
            .I3(GND_net), .O(n834_adj_2173[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_563_2 (.CI(GND_net), .I0(n598), .I1(n595), 
            .CO(n17221));
    SB_LUT4 Alpha_15__I_0_11_add_564_16_lut (.I0(GND_net), .I1(n836_adj_2182[13]), 
            .I2(n749), .I3(n17219), .O(n835[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_16 (.CI(n17219), .I0(n836_adj_2182[13]), 
            .I1(n749), .CO(n751_adj_2142));
    SB_CARRY add_1232_5 (.CI(n16903), .I0(n835_adj_2172[14]), .I1(n747_adj_2012), 
            .CO(n16904));
    SB_LUT4 add_1232_4_lut (.I0(GND_net), .I1(n834[14]), .I2(n743_adj_2096), 
            .I3(n16902), .O(Product4_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_572_2 (.CI(GND_net), .I0(n625), .I1(n622), 
            .CO(n17098));
    SB_LUT4 Alpha_15__I_0_11_add_564_15_lut (.I0(GND_net), .I1(n836_adj_2182[12]), 
            .I2(n598), .I3(n17218), .O(n835[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_15 (.CI(n17218), .I0(n836_adj_2182[12]), 
            .I1(n598), .CO(n17219));
    SB_LUT4 Alpha_15__I_0_11_add_564_14_lut (.I0(GND_net), .I1(n836_adj_2182[11]), 
            .I2(n598), .I3(n17217), .O(n835[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_14 (.CI(n17217), .I0(n836_adj_2182[11]), 
            .I1(n598), .CO(n17218));
    SB_CARRY Beta_15__I_0_add_572_2 (.CI(GND_net), .I0(n625), .I1(n622), 
            .CO(n16915));
    SB_CARRY Beta_15__I_0_add_571_3 (.CI(n16924), .I0(n843[0]), .I1(n619), 
            .CO(n16925));
    SB_LUT4 Beta_15__I_0_add_570_2_lut (.I0(GND_net), .I1(n619), .I2(n616), 
            .I3(GND_net), .O(n841[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_2 (.CI(GND_net), .I0(n619), .I1(n616), 
            .CO(n16935));
    SB_LUT4 Alpha_15__I_0_11_add_564_13_lut (.I0(GND_net), .I1(n836_adj_2182[10]), 
            .I2(n598), .I3(n17216), .O(n835[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_16_lut (.I0(GND_net), .I1(n794), .I2(n791), .I3(n17097), 
            .O(Product1_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_4_lut (.I0(GND_net), .I1(n841[1]), .I2(n613), 
            .I3(n16949), .O(n840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_3 (.CI(n16963), .I0(n840[0]), .I1(n610), 
            .CO(n16964));
    SB_CARRY Beta_15__I_0_add_568_14 (.CI(n16974), .I0(n840[11]), .I1(n610), 
            .CO(n16975));
    SB_LUT4 Beta_15__I_0_add_568_13_lut (.I0(GND_net), .I1(n840[10]), .I2(n610), 
            .I3(n16973), .O(n839[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_13 (.CI(n17216), .I0(n836_adj_2182[10]), 
            .I1(n598), .CO(n17217));
    SB_LUT4 Alpha_15__I_0_11_add_564_12_lut (.I0(GND_net), .I1(n836_adj_2182[9]), 
            .I2(n598), .I3(n17215), .O(n835[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_12 (.CI(n17215), .I0(n836_adj_2182[9]), 
            .I1(n598), .CO(n17216));
    SB_LUT4 Alpha_15__I_0_11_add_564_11_lut (.I0(GND_net), .I1(n836_adj_2182[8]), 
            .I2(n598), .I3(n17214), .O(n835[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_11 (.CI(n17214), .I0(n836_adj_2182[8]), 
            .I1(n598), .CO(n17215));
    SB_LUT4 add_1234_15_lut (.I0(GND_net), .I1(n845[14]), .I2(n787_adj_2149), 
            .I3(n17096), .O(Product1_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_13_lut (.I0(GND_net), .I1(n839[10]), .I2(n607), 
            .I3(n16988), .O(n838_adj_2170[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_566_11_lut (.I0(GND_net), .I1(n838_adj_2170[8]), 
            .I2(n604), .I3(n17001), .O(n837_adj_2171[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_564_10_lut (.I0(GND_net), .I1(n836_adj_2182[7]), 
            .I2(n598), .I3(n17213), .O(n835[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_10 (.CI(n17213), .I0(n836_adj_2182[7]), 
            .I1(n598), .CO(n17214));
    SB_CARRY Beta_15__I_0_add_565_9 (.CI(n17014), .I0(n837_adj_2171[6]), 
            .I1(n601), .CO(n17015));
    SB_CARRY add_1232_4 (.CI(n16902), .I0(n834[14]), .I1(n743_adj_2096), 
            .CO(n16903));
    SB_LUT4 Beta_15__I_0_add_565_8_lut (.I0(GND_net), .I1(n837_adj_2171[5]), 
            .I2(n601), .I3(n17013), .O(n836[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_564_9_lut (.I0(GND_net), .I1(n836_adj_2182[6]), 
            .I2(n598), .I3(n17212), .O(n835[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_9 (.CI(n17212), .I0(n836_adj_2182[6]), 
            .I1(n598), .CO(n17213));
    SB_CARRY add_1234_15 (.CI(n17096), .I0(n845[14]), .I1(n787_adj_2149), 
            .CO(n17097));
    SB_LUT4 add_1232_16_lut (.I0(GND_net), .I1(n794), .I2(n791), .I3(n16914), 
            .O(Product4_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_14_lut (.I0(GND_net), .I1(n844_adj_2181[14]), .I2(n783), 
            .I3(n17095), .O(Product1_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_564_8_lut (.I0(GND_net), .I1(n836_adj_2182[5]), 
            .I2(n598), .I3(n17211), .O(n835[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_8 (.CI(n17211), .I0(n836_adj_2182[5]), 
            .I1(n598), .CO(n17212));
    SB_CARRY add_1234_14 (.CI(n17095), .I0(n844_adj_2181[14]), .I1(n783), 
            .CO(n17096));
    SB_LUT4 Alpha_15__I_0_11_add_564_7_lut (.I0(GND_net), .I1(n836_adj_2182[4]), 
            .I2(n598), .I3(n17210), .O(n835[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_13_lut (.I0(GND_net), .I1(n843_adj_2180[14]), .I2(n779_adj_2070), 
            .I3(n17094), .O(Product1_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_7 (.CI(n17210), .I0(n836_adj_2182[4]), 
            .I1(n598), .CO(n17211));
    SB_CARRY add_1234_13 (.CI(n17094), .I0(n843_adj_2180[14]), .I1(n779_adj_2070), 
            .CO(n17095));
    SB_LUT4 add_1232_3_lut (.I0(GND_net), .I1(n833[14]), .I2(n739_adj_2006), 
            .I3(n16901), .O(Product4_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1232_15_lut (.I0(GND_net), .I1(n845[14]), .I2(n787), .I3(n16913), 
            .O(Product4_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_2_lut (.I0(GND_net), .I1(n622), .I2(n619), 
            .I3(GND_net), .O(n842[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_2 (.CI(GND_net), .I0(n622), .I1(n619), 
            .CO(n16924));
    SB_LUT4 Alpha_15__I_0_11_add_564_6_lut (.I0(GND_net), .I1(n836_adj_2182[3]), 
            .I2(n598), .I3(n17209), .O(n835[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_6 (.CI(n17209), .I0(n836_adj_2182[3]), 
            .I1(n598), .CO(n17210));
    SB_LUT4 Beta_15__I_0_add_571_12_lut (.I0(GND_net), .I1(n843[7]), .I2(n777), 
            .I3(n16933), .O(n842[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_4 (.CI(n16949), .I0(n841[1]), .I1(n613), 
            .CO(n16950));
    SB_LUT4 Beta_15__I_0_add_568_2_lut (.I0(GND_net), .I1(n613), .I2(n610), 
            .I3(GND_net), .O(n839[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_12_lut (.I0(GND_net), .I1(n842_adj_2179[14]), .I2(n775_adj_2047), 
            .I3(n17093), .O(Product1_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_2 (.CI(GND_net), .I0(n613), .I1(n610), 
            .CO(n16963));
    SB_LUT4 Alpha_15__I_0_11_add_564_5_lut (.I0(GND_net), .I1(n836_adj_2182[2]), 
            .I2(n598), .I3(n17208), .O(n835[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1234_12 (.CI(n17093), .I0(n842_adj_2179[14]), .I1(n775_adj_2047), 
            .CO(n17094));
    SB_CARRY Beta_15__I_0_add_568_13 (.CI(n16973), .I0(n840[10]), .I1(n610), 
            .CO(n16974));
    SB_CARRY Beta_15__I_0_add_567_13 (.CI(n16988), .I0(n839[10]), .I1(n607), 
            .CO(n16989));
    SB_CARRY Beta_15__I_0_add_566_11 (.CI(n17001), .I0(n838_adj_2170[8]), 
            .I1(n604), .CO(n17002));
    SB_LUT4 Beta_15__I_0_add_566_10_lut (.I0(GND_net), .I1(n838_adj_2170[7]), 
            .I2(n604), .I3(n17000), .O(n837_adj_2171[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_5 (.CI(n17208), .I0(n836_adj_2182[2]), 
            .I1(n598), .CO(n17209));
    SB_LUT4 add_1234_11_lut (.I0(GND_net), .I1(n841_adj_2178[14]), .I2(n771_adj_2032), 
            .I3(n17092), .O(Product1_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_8 (.CI(n17013), .I0(n837_adj_2171[5]), 
            .I1(n601), .CO(n17014));
    SB_LUT4 Beta_15__I_0_add_564_15_lut (.I0(GND_net), .I1(n836[12]), .I2(n598), 
            .I3(n17035), .O(n835_adj_2172[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_15 (.CI(n17035), .I0(n836[12]), .I1(n598), 
            .CO(n17036));
    SB_CARRY Beta_15__I_0_add_562_13 (.CI(n17063), .I0(n834[10]), .I1(n592), 
            .CO(n17064));
    SB_CARRY add_1234_11 (.CI(n17092), .I0(n841_adj_2178[14]), .I1(n771_adj_2032), 
            .CO(n17093));
    SB_LUT4 add_1234_10_lut (.I0(GND_net), .I1(n840_adj_2177[14]), .I2(n767), 
            .I3(n17091), .O(Product1_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_564_4_lut (.I0(GND_net), .I1(n836_adj_2182[1]), 
            .I2(n598), .I3(n17207), .O(n835[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_4 (.CI(n17207), .I0(n836_adj_2182[1]), 
            .I1(n598), .CO(n17208));
    SB_CARRY add_1234_10 (.CI(n17091), .I0(n840_adj_2177[14]), .I1(n767), 
            .CO(n17092));
    SB_LUT4 Alpha_15__I_0_11_add_564_3_lut (.I0(GND_net), .I1(n836_adj_2182[0]), 
            .I2(n598), .I3(n17206), .O(n835[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_3 (.CI(n17206), .I0(n836_adj_2182[0]), 
            .I1(n598), .CO(n17207));
    SB_LUT4 Alpha_15__I_0_11_add_564_2_lut (.I0(GND_net), .I1(n601), .I2(n598), 
            .I3(GND_net), .O(n835[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_564_2 (.CI(GND_net), .I0(n601), .I1(n598), 
            .CO(n17206));
    SB_LUT4 Alpha_15__I_0_11_add_565_16_lut (.I0(GND_net), .I1(n837[13]), 
            .I2(n753), .I3(n17204), .O(n836_adj_2182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_16 (.CI(n17204), .I0(n837[13]), .I1(n753), 
            .CO(n755_adj_2161));
    SB_LUT4 Alpha_15__I_0_11_add_565_15_lut (.I0(GND_net), .I1(n837[12]), 
            .I2(n601), .I3(n17203), .O(n836_adj_2182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_15 (.CI(n16913), .I0(n845[14]), .I1(n787), .CO(n16914));
    SB_CARRY Alpha_15__I_0_11_add_565_15 (.CI(n17203), .I0(n837[12]), .I1(n601), 
            .CO(n17204));
    SB_LUT4 Alpha_15__I_0_11_add_565_14_lut (.I0(GND_net), .I1(n837[11]), 
            .I2(n601), .I3(n17202), .O(n836_adj_2182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_14 (.CI(n17202), .I0(n837[11]), .I1(n601), 
            .CO(n17203));
    SB_LUT4 Alpha_15__I_0_11_add_565_13_lut (.I0(GND_net), .I1(n837[10]), 
            .I2(n601), .I3(n17201), .O(n836_adj_2182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_13 (.CI(n17201), .I0(n837[10]), .I1(n601), 
            .CO(n17202));
    SB_LUT4 Alpha_15__I_0_11_add_565_12_lut (.I0(GND_net), .I1(n837[9]), 
            .I2(n601), .I3(n17200), .O(n836_adj_2182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_12 (.CI(n17200), .I0(n837[9]), .I1(n601), 
            .CO(n17201));
    SB_LUT4 Alpha_15__I_0_11_add_565_11_lut (.I0(GND_net), .I1(n837[8]), 
            .I2(n601), .I3(n17199), .O(n836_adj_2182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_9_lut (.I0(GND_net), .I1(n839_adj_2174[14]), .I2(n763), 
            .I3(n17090), .O(Product1_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_12_lut (.I0(GND_net), .I1(n834[9]), .I2(n592), 
            .I3(n17062), .O(n833[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_14_lut (.I0(GND_net), .I1(n836[11]), .I2(n598), 
            .I3(n17034), .O(n835_adj_2172[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_11 (.CI(n17199), .I0(n837[8]), .I1(n601), 
            .CO(n17200));
    SB_CARRY add_1234_9 (.CI(n17090), .I0(n839_adj_2174[14]), .I1(n763), 
            .CO(n17091));
    SB_LUT4 Alpha_15__I_0_11_add_565_10_lut (.I0(GND_net), .I1(n837[7]), 
            .I2(n601), .I3(n17198), .O(n836_adj_2182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_8_lut (.I0(GND_net), .I1(n838[14]), .I2(n759_adj_2166), 
            .I3(n17089), .O(Product1_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_10 (.CI(n17198), .I0(n837[7]), .I1(n601), 
            .CO(n17199));
    SB_LUT4 Alpha_15__I_0_11_add_565_9_lut (.I0(GND_net), .I1(n837[6]), 
            .I2(n601), .I3(n17197), .O(n836_adj_2182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_3 (.CI(n16901), .I0(n833[14]), .I1(n739_adj_2006), 
            .CO(n16902));
    SB_LUT4 add_1232_14_lut (.I0(GND_net), .I1(n844[14]), .I2(n783_adj_2167), 
            .I3(n16912), .O(Product4_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1232_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1232_14 (.CI(n16912), .I0(n844[14]), .I1(n783_adj_2167), 
            .CO(n16913));
    SB_CARRY Alpha_15__I_0_11_add_565_9 (.CI(n17197), .I0(n837[6]), .I1(n601), 
            .CO(n17198));
    SB_LUT4 Beta_15__I_0_add_572_10_lut (.I0(GND_net), .I1(n844[5]), .I2(n781), 
            .I3(n16922), .O(n843[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_12 (.CI(n16933), .I0(n843[7]), .I1(n777), 
            .CO(n779));
    SB_LUT4 Beta_15__I_0_add_569_3_lut (.I0(GND_net), .I1(n841[0]), .I2(n613), 
            .I3(n16948), .O(n840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_3 (.CI(n16948), .I0(n841[0]), .I1(n613), 
            .CO(n16949));
    SB_LUT4 Alpha_15__I_0_11_add_565_8_lut (.I0(GND_net), .I1(n837[5]), 
            .I2(n601), .I3(n17196), .O(n836_adj_2182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_573_8_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n785), .I3(n17985), .O(n844_adj_2181[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_8 (.CI(n17985), .I0(n845[3]), .I1(n785), 
            .CO(n787_adj_2149));
    SB_LUT4 Alpha_15__I_0_11_add_573_7_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n625), .I3(n17984), .O(n844_adj_2181[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_7 (.CI(n17984), .I0(n845[3]), .I1(n625), 
            .CO(n17985));
    SB_LUT4 Alpha_15__I_0_11_add_573_6_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n625), .I3(n17983), .O(n844_adj_2181[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_6 (.CI(n17983), .I0(n845[3]), .I1(n625), 
            .CO(n17984));
    SB_LUT4 Alpha_15__I_0_11_add_573_5_lut (.I0(GND_net), .I1(n845[2]), 
            .I2(n625), .I3(n17982), .O(n844_adj_2181[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_5 (.CI(n17982), .I0(n845[2]), .I1(n625), 
            .CO(n17983));
    SB_LUT4 Alpha_15__I_0_11_add_573_4_lut (.I0(GND_net), .I1(n139), .I2(n625), 
            .I3(n17981), .O(n844_adj_2181[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_4 (.CI(n17981), .I0(n139), .I1(n625), 
            .CO(n17982));
    SB_LUT4 Alpha_15__I_0_11_add_573_3_lut (.I0(GND_net), .I1(n845[0]), 
            .I2(n625), .I3(n17980), .O(n844_adj_2181[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_3 (.CI(n17980), .I0(n845[0]), .I1(n625), 
            .CO(n17981));
    SB_LUT4 Alpha_15__I_0_11_add_573_2_lut (.I0(GND_net), .I1(n628), .I2(n625), 
            .I3(GND_net), .O(n844_adj_2181[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_573_2 (.CI(GND_net), .I0(n628), .I1(n625), 
            .CO(n17980));
    SB_CARRY Alpha_15__I_0_11_add_565_8 (.CI(n17196), .I0(n837[5]), .I1(n601), 
            .CO(n17197));
    SB_CARRY Beta_15__I_0_add_562_12 (.CI(n17062), .I0(n834[9]), .I1(n592), 
            .CO(n17063));
    SB_LUT4 Beta_15__I_0_add_562_11_lut (.I0(GND_net), .I1(n834[8]), .I2(n592), 
            .I3(n17061), .O(n833[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_11 (.CI(n17061), .I0(n834[8]), .I1(n592), 
            .CO(n17062));
    SB_LUT4 Alpha_15__I_0_11_add_565_7_lut (.I0(GND_net), .I1(n837[4]), 
            .I2(n601), .I3(n17195), .O(n836_adj_2182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_562_10_lut (.I0(GND_net), .I1(n834[7]), .I2(n592), 
            .I3(n17060), .O(n833[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1234_8 (.CI(n17089), .I0(n838[14]), .I1(n759_adj_2166), 
            .CO(n17090));
    SB_CARRY Alpha_15__I_0_11_add_565_7 (.CI(n17195), .I0(n837[4]), .I1(n601), 
            .CO(n17196));
    SB_LUT4 Alpha_15__I_0_11_add_565_6_lut (.I0(GND_net), .I1(n837[3]), 
            .I2(n601), .I3(n17194), .O(n836_adj_2182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_10 (.CI(n16922), .I0(n844[5]), .I1(n781), 
            .CO(n783_adj_2167));
    SB_CARRY Alpha_15__I_0_11_add_565_6 (.CI(n17194), .I0(n837[3]), .I1(n601), 
            .CO(n17195));
    SB_LUT4 Alpha_15__I_0_11_add_565_5_lut (.I0(GND_net), .I1(n837[2]), 
            .I2(n601), .I3(n17193), .O(n836_adj_2182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_5 (.CI(n17193), .I0(n837[2]), .I1(n601), 
            .CO(n17194));
    SB_LUT4 Alpha_15__I_0_11_add_565_4_lut (.I0(GND_net), .I1(n837[1]), 
            .I2(n601), .I3(n17192), .O(n836_adj_2182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_4 (.CI(n17192), .I0(n837[1]), .I1(n601), 
            .CO(n17193));
    SB_LUT4 add_1234_7_lut (.I0(GND_net), .I1(n837[14]), .I2(n755_adj_2161), 
            .I3(n17088), .O(Product1_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1234_7 (.CI(n17088), .I0(n837[14]), .I1(n755_adj_2161), 
            .CO(n17089));
    SB_LUT4 Beta_15__I_0_add_571_11_lut (.I0(GND_net), .I1(n843[7]), .I2(n619), 
            .I3(n16932), .O(n842[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_565_3_lut (.I0(GND_net), .I1(n837[0]), 
            .I2(n601), .I3(n17191), .O(n836_adj_2182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_565_3 (.CI(n17191), .I0(n837[0]), .I1(n601), 
            .CO(n17192));
    SB_LUT4 Alpha_15__I_0_11_add_565_2_lut (.I0(GND_net), .I1(n604), .I2(n601), 
            .I3(GND_net), .O(n836_adj_2182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_10 (.CI(n17060), .I0(n834[7]), .I1(n592), 
            .CO(n17061));
    SB_CARRY Alpha_15__I_0_11_add_565_2 (.CI(GND_net), .I0(n604), .I1(n601), 
            .CO(n17191));
    SB_LUT4 Alpha_15__I_0_11_add_566_16_lut (.I0(GND_net), .I1(n838[13]), 
            .I2(n757), .I3(n17189), .O(n837[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1234_6_lut (.I0(GND_net), .I1(n836_adj_2182[14]), .I2(n751_adj_2142), 
            .I3(n17087), .O(Product1_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1234_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_2_lut (.I0(GND_net), .I1(n616), .I2(n613), 
            .I3(GND_net), .O(n840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_16 (.CI(n17189), .I0(n838[13]), .I1(n757), 
            .CO(n759_adj_2166));
    SB_LUT4 Alpha_15__I_0_11_add_566_15_lut (.I0(GND_net), .I1(n838[12]), 
            .I2(n604), .I3(n17188), .O(n837[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_15 (.CI(n17188), .I0(n838[12]), .I1(n604), 
            .CO(n17189));
    SB_CARRY Beta_15__I_0_add_569_2 (.CI(GND_net), .I0(n616), .I1(n613), 
            .CO(n16948));
    SB_LUT4 Beta_15__I_0_add_562_9_lut (.I0(GND_net), .I1(n834[6]), .I2(n592), 
            .I3(n17059), .O(n833[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_add_566_14_lut (.I0(GND_net), .I1(n838[11]), 
            .I2(n604), .I3(n17187), .O(n837[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_14 (.CI(n17187), .I0(n838[11]), .I1(n604), 
            .CO(n17188));
    SB_LUT4 Alpha_15__I_0_11_add_566_13_lut (.I0(GND_net), .I1(n838[10]), 
            .I2(n604), .I3(n17186), .O(n837[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_13 (.CI(n17186), .I0(n838[10]), .I1(n604), 
            .CO(n17187));
    SB_LUT4 Alpha_15__I_0_11_add_566_12_lut (.I0(GND_net), .I1(n838[9]), 
            .I2(n604), .I3(n17185), .O(n837[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_11_add_566_12 (.CI(n17185), .I0(n838[9]), .I1(n604), 
            .CO(n17186));
    SB_LUT4 sub_65_add_2_29_lut (.I0(GND_net), .I1(Product4_mul_temp[29]), 
            .I2(VCC_net), .I3(n15774), .O(\qCurrent[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_65_add_2_28_lut (.I0(GND_net), .I1(Product4_mul_temp[28]), 
            .I2(VCC_net), .I3(n15773), .O(\qCurrent[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_28 (.CI(n15773), .I0(Product4_mul_temp[28]), .I1(VCC_net), 
            .CO(n15774));
    SB_LUT4 sub_65_add_2_27_lut (.I0(GND_net), .I1(Product4_mul_temp[27]), 
            .I2(VCC_net), .I3(n15772), .O(\qCurrent[29] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_27 (.CI(n15772), .I0(Product4_mul_temp[27]), .I1(VCC_net), 
            .CO(n15773));
    SB_LUT4 sub_65_add_2_26_lut (.I0(GND_net), .I1(Product4_mul_temp[26]), 
            .I2(VCC_net), .I3(n15771), .O(\qCurrent[28] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_26 (.CI(n15771), .I0(Product4_mul_temp[26]), .I1(VCC_net), 
            .CO(n15772));
    SB_LUT4 sub_65_add_2_25_lut (.I0(GND_net), .I1(Product4_mul_temp[25]), 
            .I2(VCC_net), .I3(n15770), .O(\qCurrent[27] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_25 (.CI(n15770), .I0(Product4_mul_temp[25]), .I1(VCC_net), 
            .CO(n15771));
    SB_LUT4 sub_65_add_2_24_lut (.I0(GND_net), .I1(Product4_mul_temp[24]), 
            .I2(VCC_net), .I3(n15769), .O(\qCurrent[26] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_24 (.CI(n15769), .I0(Product4_mul_temp[24]), .I1(VCC_net), 
            .CO(n15770));
    SB_LUT4 sub_65_add_2_23_lut (.I0(GND_net), .I1(Product4_mul_temp[23]), 
            .I2(VCC_net), .I3(n15768), .O(\qCurrent[25] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_23 (.CI(n15768), .I0(Product4_mul_temp[23]), .I1(VCC_net), 
            .CO(n15769));
    SB_LUT4 sub_65_add_2_22_lut (.I0(GND_net), .I1(Product4_mul_temp[22]), 
            .I2(VCC_net), .I3(n15767), .O(\qCurrent[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_22 (.CI(n15767), .I0(Product4_mul_temp[22]), .I1(VCC_net), 
            .CO(n15768));
    SB_LUT4 sub_65_add_2_21_lut (.I0(GND_net), .I1(Product4_mul_temp[21]), 
            .I2(VCC_net), .I3(n15766), .O(\qCurrent[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_21 (.CI(n15766), .I0(Product4_mul_temp[21]), .I1(VCC_net), 
            .CO(n15767));
    SB_LUT4 sub_65_add_2_20_lut (.I0(GND_net), .I1(Product4_mul_temp[20]), 
            .I2(VCC_net), .I3(n15765), .O(\qCurrent[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_20 (.CI(n15765), .I0(Product4_mul_temp[20]), .I1(VCC_net), 
            .CO(n15766));
    SB_LUT4 sub_65_add_2_19_lut (.I0(GND_net), .I1(Product4_mul_temp[19]), 
            .I2(VCC_net), .I3(n15764), .O(\qCurrent[21] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_i498_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i498_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY sub_65_add_2_19 (.CI(n15764), .I0(Product4_mul_temp[19]), .I1(VCC_net), 
            .CO(n15765));
    SB_LUT4 sub_65_add_2_18_lut (.I0(GND_net), .I1(Product4_mul_temp[18]), 
            .I2(VCC_net), .I3(n15763), .O(\qCurrent[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_18 (.CI(n15763), .I0(Product4_mul_temp[18]), .I1(VCC_net), 
            .CO(n15764));
    SB_LUT4 sub_65_add_2_17_lut (.I0(GND_net), .I1(Product4_mul_temp[17]), 
            .I2(VCC_net), .I3(n15762), .O(\qCurrent[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_17 (.CI(n15762), .I0(Product4_mul_temp[17]), .I1(VCC_net), 
            .CO(n15763));
    SB_LUT4 sub_65_add_2_16_lut (.I0(GND_net), .I1(Product4_mul_temp[16]), 
            .I2(VCC_net), .I3(n15761), .O(\qCurrent[18] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_16 (.CI(n15761), .I0(Product4_mul_temp[16]), .I1(VCC_net), 
            .CO(n15762));
    SB_LUT4 sub_65_add_2_15_lut (.I0(GND_net), .I1(Product4_mul_temp[15]), 
            .I2(VCC_net), .I3(n15760), .O(\qCurrent[17] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_15 (.CI(n15760), .I0(Product4_mul_temp[15]), .I1(VCC_net), 
            .CO(n15761));
    SB_LUT4 sub_65_add_2_14_lut (.I0(GND_net), .I1(Product4_mul_temp[14]), 
            .I2(VCC_net), .I3(n15759), .O(\qCurrent[16] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_i12_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n604));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Alpha_15__I_0_11_i22_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n619));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_65_add_2_14 (.CI(n15759), .I0(Product4_mul_temp[14]), .I1(VCC_net), 
            .CO(n15760));
    SB_LUT4 sub_65_add_2_13_lut (.I0(GND_net), .I1(Product4_mul_temp[13]), 
            .I2(VCC_net), .I3(n15758), .O(\qCurrent[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_13 (.CI(n15758), .I0(Product4_mul_temp[13]), .I1(VCC_net), 
            .CO(n15759));
    SB_LUT4 sub_65_add_2_12_lut (.I0(GND_net), .I1(Product4_mul_temp[12]), 
            .I2(VCC_net), .I3(n15757), .O(\qCurrent[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_12 (.CI(n15757), .I0(Product4_mul_temp[12]), .I1(VCC_net), 
            .CO(n15758));
    SB_LUT4 sub_65_add_2_11_lut (.I0(GND_net), .I1(Product4_mul_temp[11]), 
            .I2(VCC_net), .I3(n15756), .O(\qCurrent[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_11 (.CI(n15756), .I0(Product4_mul_temp[11]), .I1(VCC_net), 
            .CO(n15757));
    SB_LUT4 sub_65_add_2_10_lut (.I0(GND_net), .I1(Product4_mul_temp[10]), 
            .I2(VCC_net), .I3(n15755), .O(\qCurrent[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_10 (.CI(n15755), .I0(Product4_mul_temp[10]), .I1(VCC_net), 
            .CO(n15756));
    SB_LUT4 sub_65_add_2_9_lut (.I0(GND_net), .I1(Product4_mul_temp[9]), 
            .I2(VCC_net), .I3(n15754), .O(\qCurrent[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_9 (.CI(n15754), .I0(Product4_mul_temp[9]), .I1(VCC_net), 
            .CO(n15755));
    SB_LUT4 sub_65_add_2_8_lut (.I0(GND_net), .I1(Product4_mul_temp[8]), 
            .I2(VCC_net), .I3(n15753), .O(\qCurrent[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_8 (.CI(n15753), .I0(Product4_mul_temp[8]), .I1(VCC_net), 
            .CO(n15754));
    SB_LUT4 sub_65_add_2_7_lut (.I0(GND_net), .I1(Product4_mul_temp[7]), 
            .I2(VCC_net), .I3(n15752), .O(\qCurrent[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_7 (.CI(n15752), .I0(Product4_mul_temp[7]), .I1(VCC_net), 
            .CO(n15753));
    SB_LUT4 sub_65_add_2_6_lut (.I0(GND_net), .I1(Product4_mul_temp[6]), 
            .I2(VCC_net), .I3(n15751), .O(\qCurrent[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_6 (.CI(n15751), .I0(Product4_mul_temp[6]), .I1(VCC_net), 
            .CO(n15752));
    SB_LUT4 sub_65_add_2_5_lut (.I0(GND_net), .I1(Product4_mul_temp[5]), 
            .I2(VCC_net), .I3(n15750), .O(\qCurrent[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_5 (.CI(n15750), .I0(Product4_mul_temp[5]), .I1(VCC_net), 
            .CO(n15751));
    SB_LUT4 sub_65_add_2_4_lut (.I0(GND_net), .I1(Product4_mul_temp[4]), 
            .I2(VCC_net), .I3(n15749), .O(\qCurrent[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_4 (.CI(n15749), .I0(Product4_mul_temp[4]), .I1(VCC_net), 
            .CO(n15750));
    SB_LUT4 sub_65_add_2_3_lut (.I0(GND_net), .I1(Product4_mul_temp[3]), 
            .I2(VCC_net), .I3(n15748), .O(\qCurrent[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_3 (.CI(n15748), .I0(Product4_mul_temp[3]), .I1(VCC_net), 
            .CO(n15749));
    SB_LUT4 sub_65_add_2_2_lut (.I0(GND_net), .I1(Product4_mul_temp[2]), 
            .I2(\Amp25_out1[14] ), .I3(VCC_net), .O(\qCurrent[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_65_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_65_add_2_2 (.CI(VCC_net), .I0(Product4_mul_temp[2]), .I1(\Amp25_out1[14] ), 
            .CO(n15748));
    SB_LUT4 Beta_15__I_0_i528_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n777));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i528_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Beta_15__I_0_i516_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i516_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY Beta_15__I_0_add_562_9 (.CI(n17059), .I0(n834[6]), .I1(n592), 
            .CO(n17060));
    SB_CARRY add_1234_6 (.CI(n17087), .I0(n836_adj_2182[14]), .I1(n751_adj_2142), 
            .CO(n17088));
    SB_LUT4 Alpha_15__I_0_11_add_566_11_lut (.I0(GND_net), .I1(n838[8]), 
            .I2(n604), .I3(n17184), .O(n837[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_11_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_11_i18_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n613));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Alpha_15__I_0_11_i8_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n598));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Beta_15__I_0_i513_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n757));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i513_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Beta_15__I_0_i510_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n753));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i510_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_4_lut (.I0(n142), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_out1_1[13]), 
            .I3(n26), .O(n845[14]));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h4c26;
    SB_LUT4 Beta_15__I_0_i525_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n773));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i525_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Alpha_15__I_0_11_i14_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n607));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Beta_15__I_0_i522_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n769));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(66[30:52])
    defparam Beta_15__I_0_i522_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Alpha_15__I_0_11_i16_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n610));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(n142), .I1(\Product_mul_temp[26] ), 
            .I2(Look_Up_Table_out1_1[13]), .I3(n4), .O(n12));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 Alpha_15__I_0_11_i4_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n592));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam Alpha_15__I_0_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_3_lut_4_lut (.I0(n142), .I1(\Product_mul_temp[26] ), 
            .I2(Look_Up_Table_out1_1[13]), .I3(n4), .O(n6));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_3_lut_3_lut_4_lut.LUT_INIT = 16'haa80;
    SB_LUT4 i1_3_lut_4_lut (.I0(n4), .I1(n142), .I2(\Product_mul_temp[26] ), 
            .I3(Look_Up_Table_out1_1[13]), .O(n845[3]));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hd444;
    SB_LUT4 i2_3_lut_4_lut (.I0(n4), .I1(\Product_mul_temp[26] ), .I2(Look_Up_Table_out1_1[13]), 
            .I3(n142), .O(n845[2]));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 i1_3_lut_4_lut_adj_308 (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(n6), .I3(n12), .O(n14));   // ../../hdlcoderFocCurrentFixptHdl/Park_Transform.v(50[30:53])
    defparam i1_3_lut_4_lut_adj_308.LUT_INIT = 16'hf8f0;
    VCC i1 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module Inverse_Park_Transform
//

module Inverse_Park_Transform (\qVoltage[6] , Look_Up_Table_out1_1, GND_net, 
            \dVoltage[11] , \qVoltage[7] , n610, \Product_mul_temp[26] , 
            \qVoltage[9] , \Product2_mul_temp[2] , n86, \dVoltage[6] , 
            \qVoltage[10] , n576, n414, n267, n218, \qVoltage[13] , 
            \qVoltage[14] , \qVoltage[12] , n236, n120, \qVoltage[3] , 
            \dVoltage[10] , \qVoltage[4] , \Product3_mul_temp[2] , n26, 
            n71, n138, n44, n89, \betaVoltage[15] , n209, \betaVoltage[14] , 
            n19681, n19684, n769, n685, n587, n631, \betaVoltage[13] , 
            n264, n114, n613, n417, \betaVoltage[12] , \qVoltage[8] , 
            n270, n221, n123, n29, n74, n773, n616, n420, \betaVoltage[11] , 
            n273, n224, n126, n32, n77, n777, n619, n587_adj_203, 
            n489, n391, n342, \dVoltage[15] , n233, n86_adj_204, 
            n423, n276, n227, n538, n685_adj_205, n587_adj_206, 
            n489_adj_207, n391_adj_208, n342_adj_209, n244, n129, 
            n35, n80, n781, n489_adj_210, n622, n215, n11, n56, 
            n749, \qVoltage[15] , n102, n592, n393, n391_adj_211, 
            n435, n255, n342_adj_212, n737, n20, n65, n111, n405, 
            n206, n737_adj_213, n598, n399, n8, n53, \dVoltage[9] , 
            n589, n540, n393_adj_214, n246, n99, n19351, n50, 
            n741, n592_adj_215, n543, n396, n249, n102_adj_216, 
            n8_adj_217, n53_adj_218, n745, n595, n546, n399_adj_219, 
            n252, n105, n11_adj_220, n56_adj_221, n749_adj_222, n598_adj_223, 
            n549, n402, n255_adj_224, n108, n14, n59, n753, n601, 
            n552, n405_adj_225, n258, n111_adj_226, n17, n62, n757, 
            n604, n555, n408, n261, n114_adj_227, n20_adj_228, n65_adj_229, 
            n761, n607, n558, n411, n264_adj_230, n117, n23, n68, 
            n765, n610_adj_231, n561, n414_adj_232, n267_adj_233, 
            n761_adj_234, n120_adj_235, n26_adj_236, n71_adj_237, n769_adj_238, 
            n613_adj_239, n564, n417_adj_240, n17_adj_241, n62_adj_242, 
            n601_adj_243, n244_adj_244, n288, n195, n239, alphaVoltage, 
            n408_adj_245, n108_adj_246, n402_adj_247, n270_adj_248, 
            n745_adj_249, n141, n246_adj_250, n123_adj_251, n117_adj_252, 
            n757_adj_253, n23_adj_254, n68_adj_255, n252_adj_256, n396_adj_257, 
            n92, n197, n29_adj_258, n74_adj_259, n773_adj_260, n616_adj_261, 
            n567, \dVoltage[5] , n420_adj_262, n273_adj_263, n126_adj_264, 
            n32_adj_265, n77_adj_266, n777_adj_267, n619_adj_268, n570, 
            n423_adj_269, n276_adj_270, n129_adj_271, n35_adj_272, n80_adj_273, 
            n781_adj_274, n622_adj_275, n573, n426, n279, n132, 
            n38, n83, n785, n625, n576_adj_276, n589_adj_277, n429, 
            n282, n135, n41, n86_adj_278, n789, n628, n579, n432, 
            n285, n138_adj_279, n44_adj_280, n89_adj_281, n19604, 
            n685_adj_282, n587_adj_283, n631_adj_284, n538_adj_285, 
            n582, n489_adj_286, n391_adj_287, n435_adj_288, n342_adj_289, 
            n244_adj_290, n288_adj_291, n195_adj_292, n141_adj_293, 
            n92_adj_294, \betaVoltage[10] , n203, n99_adj_295, \dVoltage[14] , 
            \dVoltage[7] , \dVoltage[3] , \dVoltage[13] , \betaVoltage[9] , 
            n19576, n50_adj_296, \betaVoltage[8] , n261_adj_297, n19702, 
            n595_adj_298, n249_adj_299, n741_adj_300, Out_31__N_333, 
            \preSatVoltage[10] , Out_31__N_332, \qVoltage[2] , \qVoltage[5] , 
            \dVoltage[8] , n426_adj_301, n258_adj_302, \preSatVoltage[13] , 
            \preSatVoltage[12] , \preSatVoltage[19] , \preSatVoltage[22] , 
            \preSatVoltage[23] , n19352, Out_31__N_333_adj_303, \preSatVoltage[10]_adj_304 , 
            Out_31__N_332_adj_305, \dVoltage[2] , n411_adj_306, n14_adj_307, 
            n59_adj_308, n200, n753_adj_309, n105_adj_310, n765_adj_311, 
            n607_adj_312, n212, n604_adj_313, \betaVoltage[7] , \betaVoltage[6] , 
            n279_adj_314, n230, n132_adj_315, n38_adj_316, n83_adj_317, 
            n785_adj_318, \dVoltage[12] , \betaVoltage[5] , n625_adj_319, 
            \betaVoltage[4] , \betaVoltage[3] , \betaVoltage[2] , \Gain1_mul_temp[2] , 
            \Gain1_mul_temp[1] , n429_adj_320, \preSatVoltage[23]_adj_321 , 
            \preSatVoltage[19]_adj_322 , \preSatVoltage[12]_adj_323 , n282_adj_324, 
            n233_adj_325, n135_adj_326, n41_adj_327, n86_adj_328, n789_adj_329, 
            n628_adj_330, n432_adj_331, n285_adj_332) /* synthesis syn_module_defined=1 */ ;
    input \qVoltage[6] ;
    input [15:0]Look_Up_Table_out1_1;
    input GND_net;
    input \dVoltage[11] ;
    input \qVoltage[7] ;
    input n610;
    input \Product_mul_temp[26] ;
    input \qVoltage[9] ;
    input \Product2_mul_temp[2] ;
    input n86;
    input \dVoltage[6] ;
    input \qVoltage[10] ;
    input n576;
    input n414;
    input n267;
    input n218;
    input \qVoltage[13] ;
    input \qVoltage[14] ;
    input \qVoltage[12] ;
    input n236;
    input n120;
    input \qVoltage[3] ;
    input \dVoltage[10] ;
    input \qVoltage[4] ;
    input \Product3_mul_temp[2] ;
    input n26;
    input n71;
    input n138;
    input n44;
    input n89;
    output \betaVoltage[15] ;
    input n209;
    output \betaVoltage[14] ;
    input n19681;
    input n19684;
    input n769;
    input n685;
    input n587;
    input n631;
    output \betaVoltage[13] ;
    input n264;
    input n114;
    input n613;
    input n417;
    output \betaVoltage[12] ;
    input \qVoltage[8] ;
    input n270;
    input n221;
    input n123;
    input n29;
    input n74;
    input n773;
    input n616;
    input n420;
    output \betaVoltage[11] ;
    input n273;
    input n224;
    input n126;
    input n32;
    input n77;
    input n777;
    input n619;
    input n587_adj_203;
    input n489;
    input n391;
    input n342;
    input \dVoltage[15] ;
    input n233;
    input n86_adj_204;
    input n423;
    input n276;
    input n227;
    input n538;
    input n685_adj_205;
    input n587_adj_206;
    input n489_adj_207;
    input n391_adj_208;
    input n342_adj_209;
    input n244;
    input n129;
    input n35;
    input n80;
    input n781;
    input n489_adj_210;
    input n622;
    input n215;
    input n11;
    input n56;
    input n749;
    input \qVoltage[15] ;
    input n102;
    input n592;
    input n393;
    input n391_adj_211;
    input n435;
    input n255;
    input n342_adj_212;
    input n737;
    input n20;
    input n65;
    input n111;
    input n405;
    input n206;
    input n737_adj_213;
    input n598;
    input n399;
    input n8;
    input n53;
    input \dVoltage[9] ;
    input n589;
    input n540;
    input n393_adj_214;
    input n246;
    input n99;
    input n19351;
    input n50;
    input n741;
    input n592_adj_215;
    input n543;
    input n396;
    input n249;
    input n102_adj_216;
    input n8_adj_217;
    input n53_adj_218;
    input n745;
    input n595;
    input n546;
    input n399_adj_219;
    input n252;
    input n105;
    input n11_adj_220;
    input n56_adj_221;
    input n749_adj_222;
    input n598_adj_223;
    input n549;
    input n402;
    input n255_adj_224;
    input n108;
    input n14;
    input n59;
    input n753;
    input n601;
    input n552;
    input n405_adj_225;
    input n258;
    input n111_adj_226;
    input n17;
    input n62;
    input n757;
    input n604;
    input n555;
    input n408;
    input n261;
    input n114_adj_227;
    input n20_adj_228;
    input n65_adj_229;
    input n761;
    input n607;
    input n558;
    input n411;
    input n264_adj_230;
    input n117;
    input n23;
    input n68;
    input n765;
    input n610_adj_231;
    input n561;
    input n414_adj_232;
    input n267_adj_233;
    input n761_adj_234;
    input n120_adj_235;
    input n26_adj_236;
    input n71_adj_237;
    input n769_adj_238;
    input n613_adj_239;
    input n564;
    input n417_adj_240;
    input n17_adj_241;
    input n62_adj_242;
    input n601_adj_243;
    input n244_adj_244;
    input n288;
    input n195;
    input n239;
    output [15:0]alphaVoltage;
    input n408_adj_245;
    input n108_adj_246;
    input n402_adj_247;
    input n270_adj_248;
    input n745_adj_249;
    input n141;
    input n246_adj_250;
    input n123_adj_251;
    input n117_adj_252;
    input n757_adj_253;
    input n23_adj_254;
    input n68_adj_255;
    input n252_adj_256;
    input n396_adj_257;
    input n92;
    input n197;
    input n29_adj_258;
    input n74_adj_259;
    input n773_adj_260;
    input n616_adj_261;
    input n567;
    input \dVoltage[5] ;
    input n420_adj_262;
    input n273_adj_263;
    input n126_adj_264;
    input n32_adj_265;
    input n77_adj_266;
    input n777_adj_267;
    input n619_adj_268;
    input n570;
    input n423_adj_269;
    input n276_adj_270;
    input n129_adj_271;
    input n35_adj_272;
    input n80_adj_273;
    input n781_adj_274;
    input n622_adj_275;
    input n573;
    input n426;
    input n279;
    input n132;
    input n38;
    input n83;
    input n785;
    input n625;
    input n576_adj_276;
    input n589_adj_277;
    input n429;
    input n282;
    input n135;
    input n41;
    input n86_adj_278;
    input n789;
    input n628;
    input n579;
    input n432;
    input n285;
    input n138_adj_279;
    input n44_adj_280;
    input n89_adj_281;
    input n19604;
    input n685_adj_282;
    input n587_adj_283;
    input n631_adj_284;
    input n538_adj_285;
    input n582;
    input n489_adj_286;
    input n391_adj_287;
    input n435_adj_288;
    input n342_adj_289;
    input n244_adj_290;
    input n288_adj_291;
    input n195_adj_292;
    input n141_adj_293;
    input n92_adj_294;
    output \betaVoltage[10] ;
    input n203;
    input n99_adj_295;
    input \dVoltage[14] ;
    input \dVoltage[7] ;
    input \dVoltage[3] ;
    input \dVoltage[13] ;
    output \betaVoltage[9] ;
    input n19576;
    input n50_adj_296;
    output \betaVoltage[8] ;
    input n261_adj_297;
    input n19702;
    input n595_adj_298;
    input n249_adj_299;
    input n741_adj_300;
    input Out_31__N_333;
    input \preSatVoltage[10] ;
    input Out_31__N_332;
    input \qVoltage[2] ;
    input \qVoltage[5] ;
    input \dVoltage[8] ;
    input n426_adj_301;
    input n258_adj_302;
    input \preSatVoltage[13] ;
    input \preSatVoltage[12] ;
    input \preSatVoltage[19] ;
    input \preSatVoltage[22] ;
    input \preSatVoltage[23] ;
    input n19352;
    input Out_31__N_333_adj_303;
    input \preSatVoltage[10]_adj_304 ;
    input Out_31__N_332_adj_305;
    input \dVoltage[2] ;
    input n411_adj_306;
    input n14_adj_307;
    input n59_adj_308;
    input n200;
    input n753_adj_309;
    input n105_adj_310;
    input n765_adj_311;
    input n607_adj_312;
    input n212;
    input n604_adj_313;
    output \betaVoltage[7] ;
    output \betaVoltage[6] ;
    input n279_adj_314;
    input n230;
    input n132_adj_315;
    input n38_adj_316;
    input n83_adj_317;
    input n785_adj_318;
    input \dVoltage[12] ;
    output \betaVoltage[5] ;
    input n625_adj_319;
    output \betaVoltage[4] ;
    output \betaVoltage[3] ;
    output \betaVoltage[2] ;
    output \Gain1_mul_temp[2] ;
    output \Gain1_mul_temp[1] ;
    input n429_adj_320;
    input \preSatVoltage[23]_adj_321 ;
    input \preSatVoltage[19]_adj_322 ;
    input \preSatVoltage[12]_adj_323 ;
    input n282_adj_324;
    input n233_adj_325;
    input n135_adj_326;
    input n41_adj_327;
    input n86_adj_328;
    input n789_adj_329;
    input n628_adj_330;
    input n432_adj_331;
    input n285_adj_332;
    
    
    wire n310;
    wire [14:0]n842;
    wire [14:0]n843;
    
    wire n331, n16545, n546_c, n16546, n359, n282_c, n16544, n233_c, 
        n16543, n184, n16542;
    wire [14:0]n839;
    wire [14:0]n840;
    
    wire n16588, n16790;
    wire [14:0]n840_adj_1950;
    
    wire n16791, n16552, n674, n16553, n135_c, n16541, n380, n457, 
        n17676;
    wire [31:0]Product3_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(46[22:39])
    wire [31:0]Product4_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(48[22:39])
    
    wire n17677;
    wire [14:0]n844;
    
    wire n793, n16539, n783, n723, n16538;
    wire [14:0]n839_adj_1951;
    
    wire n561_c, n16789, n17675, n16537, n17674, n625_c, n16536, 
        n304, n506, n16535, n527, n16534, n16589, n512, n16788, 
        n463, n16787, n16786, n365, n16785, n316, n16784, n16783, 
        n16782, n16655;
    wire [14:0]n836;
    
    wire n16656, n653, n702, n16692;
    wire [14:0]n846;
    
    wire n16693, n169, n16781, n16587;
    wire [14:0]n835;
    
    wire n16654, n17673, n16780, n160, n478, n16653, n491, n17672, 
        n209_c, n307, n356, n17671, n17670, n17669, n16533;
    wire [14:0]n845;
    
    wire n187, n16691;
    wire [31:0]Product2_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(40[22:39])
    
    wire n16661, n16556, n16690, n16662, n17696, n16827;
    wire [14:0]n837;
    
    wire n16828, n16586, n17695, n16689;
    wire [14:0]n841;
    
    wire n16778, n16554, n779, n429_c, n16532, n454, n16531, n503, 
        n771, n729, n16688;
    wire [14:0]n841_adj_1952;
    
    wire n16584, n636, n680, n16687, n771_adj_1019, n711, n16777, 
        n16686, n662, n16776, n17694, n503_adj_1020, n16799, n313, 
        n16800;
    wire [14:0]n838;
    
    wire n16798, n16810, n16792, n708, n16793, n16530, n16583, 
        n650;
    wire [14:0]n838_adj_1953;
    
    wire n16612, n16613, n16614, n699, n16611, n16582, n16610, 
        n16609, n16608, n16652, n16775, n564_c, n16774, n157, 
        n515, n16773, n16651, n466, n16772, n16771, n16650, n206_c, 
        n368, n16770, n16649, n319, n16769, n16581, n304_adj_1031, 
        n16607, n16606, n353, n16605, n451, n17693, n500, n16604, 
        n16603, n16648, n16768, n16767, n172, n16766, n16647, 
        n16765, n16646, n647, n696;
    wire [14:0]n842_adj_1954;
    
    wire n16763, n775, n714, n16762;
    wire [14:0]n837_adj_1955;
    
    wire n16644, n665, n16761, n16760, n567_c, n16759, n518, n16758, 
        n469, n16757, n16756, n154, n16577, n16578, n16579, n16580, 
        n203_c, n16602, n17692, n16601, n301, n350, n16574, n16575, 
        n16576, n448, n497, n755, n371, n16755, n16643, n322, 
        n16754, n16642, n16753, n16752, n175, n16751, n16750, 
        n16571, n16572, n16573, n644, n16599, n767, n693, n16598, 
        n16567, n16568, n16569, n775_adj_1064, n16641, n16640;
    wire [14:0]n843_adj_1956;
    
    wire n16748, n779_adj_1067, n16639, n717, n16747, n668, n16746, 
        n16745, n16529, n16528, n570_c, n16744, n16638, n16637, 
        n16527, n16526;
    wire [14:0]n845_adj_1957;
    
    wire n16524, n787, n16523, n16522, n151, n16521, n16520, n16519, 
        n200_c, n298, n347, n16518, n445, n494, n16517, n16516, 
        n16515, n16514, n16513, n16512, n16511, n16636;
    wire [14:0]n846_adj_1958;
    
    wire n16509, n791, n641, n690, n16508, n16507, n16506, n16505, 
        n16504, n16503, n16502, n16501, n16500, n16499, n16635, 
        n16498, n16497, n16496, n19680, n16495, n685_adj_1082, n16494, 
        n636_adj_1083, n16493, n16492, n538_c, n16491, n16490, n440, 
        n16489, n16488, n16487, n16634, n293, n16486, n16633, 
        n244_c, n16485, n195_c, n16484, n146, n16483, n97, n16482, 
        n48;
    wire [31:0]Product1_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(38[22:39])
    
    wire n791_adj_1086, n16481, n787_adj_1088, n16480;
    wire [14:0]n844_adj_1959;
    
    wire n783_adj_1090, n16479, n16478, n16477, n16476, n767_adj_1092, 
        n16475, n763, n16474, n759, n16473, n755_adj_1094, n16472;
    wire [14:0]n836_adj_1960;
    
    wire n751, n16471;
    wire [14:0]n835_adj_1961;
    
    wire n747, n16470, n521, n16743;
    wire [14:0]n834;
    
    wire n743, n16469;
    wire [14:0]n833;
    
    wire n739, n16468, n16467;
    wire [14:0]n832;
    wire [14:0]n834_adj_1962;
    wire [14:0]n835_adj_1963;
    
    wire n793_adj_1098, n16465, n747_adj_1099, n723_adj_1100, n16464;
    wire [14:0]n833_adj_1964;
    
    wire n674_adj_1101, n16463, n625_adj_1102, n16462, n576_adj_1104, 
        n16461, n527_adj_1106, n16460, n478_adj_1108, n16459, n429_adj_1110, 
        n16458, n380_adj_1112, n16457, n331_adj_1114, n16456, n282_adj_1116, 
        n16455, n16454, n184_adj_1120, n16453, n16632, n135_adj_1123, 
        n16452;
    wire [14:0]n836_adj_1965;
    
    wire n16450, n751_adj_1127, n16449, n16448, n16447, n472, n16742, 
        n16446, n16445, n16444, n16443, n16442, n16441, n16440, 
        n16439, n16438, n16437;
    wire [14:0]n837_adj_1966;
    
    wire n16435, n755_adj_1144, n16434, n16433, n16432, n16431, 
        n16430, n16429, n16428, n16427, n16426, n16425, n16424, 
        n16423, n16422;
    wire [14:0]n838_adj_1967;
    
    wire n16420, n759_adj_1158, n16419, n16418, n16417, n16416, 
        n16415, n16414, n16413, n16412, n16411, n16410, n16409, 
        n16631, n16408, n16407;
    wire [14:0]n839_adj_1968;
    
    wire n16405, n763_adj_1175, n16404, n16403, n16402, n16401, 
        n16400, n16399, n16398, n16397, n16396, n16395, n16394, 
        n16393, n16392;
    wire [14:0]n840_adj_1969;
    
    wire n16390, n767_adj_1191, n16389, n16388, n16387, n16386, 
        n16385, n16384, n16383, n16382, n16381, n16380, n16379, 
        n16378, n16377;
    wire [14:0]n841_adj_1970;
    
    wire n16375, n771_adj_1207, n16374, n16373, n16372, n16371, 
        n16370, n16369, n16368, n16367, n16741, n16366, n16365, 
        n16364, n16363, n16362;
    wire [14:0]n842_adj_1971;
    
    wire n16360, n775_adj_1224, n16359, n16358, n374, n16740, n16357, 
        n16356, n16355, n16354, n16353, n16352, n16351, n16350, 
        n16349, n16348, n16347;
    wire [14:0]n843_adj_1972;
    
    wire n16345, n779_adj_1241, n16344, n16343, n16342, n16341, 
        n16340, n16339, n16338, n16337, n16336, n16335, n16334, 
        n16333, n16332;
    wire [14:0]n844_adj_1973;
    
    wire n16330, n783_adj_1257, n16329, n16328, n16327, n16326, 
        n16325, n16324, n16323, n16322, n16321, n16320, n16319, 
        n16318, n16317;
    wire [14:0]n845_adj_1974;
    
    wire n16315, n787_adj_1273, n16314, n16313, n16312, n16311, 
        n16310, n16309, n16308, n16307, n16306, n16305, n16304, 
        n16303, n16302;
    wire [14:0]n846_adj_1975;
    
    wire n16300, n791_adj_1289, n16299, n16298, n325, n16739, n16297, 
        n16296, n16295, n16294, n16293, n16292, n16291, n16290, 
        n16738, n16289, n16288, n16287, n16737, n19585, n16286, 
        n16597, n582_c, n16685, n16285, n636_adj_1310, n16284, n16283, 
        n538_adj_1312, n16282, n148, n16281, n197_c, n440_adj_1314, 
        n16280, n16279, n16278, n293_adj_1317, n16277, n178, n16736, 
        n16276, n195_adj_1320, n16275, n146_adj_1321, n16274, n97_adj_1322, 
        n16273, n16629, n16735, n48_adj_1326, n16272, n16271, n759_adj_1327, 
        n295, n16270, n16269, n16733, n16268, n344, n442, n491_adj_1330, 
        n16267, n16266, n763_adj_1331, n16265, n16264, n638, n295_adj_1333, 
        n16263, n751_adj_1334, n16262, n720, n16732, n747_adj_1337, 
        n16261, n533, n16684, n16596, n440_adj_1341, n484, n16683, 
        n16566;
    wire [14:0]n834_adj_1976;
    
    wire n9636, n16260, n671, n16731, n16628, n16730;
    wire [14:0]n833_adj_1977;
    
    wire n9213, n16259, n659, n16797, n16855, n16853, n16258, 
        n16863, n497_adj_1351, n16864, n16870;
    wire [14:0]n832_adj_1978;
    
    wire n16881, n641_adj_1353, n16882, n16257, n16256, n16255, 
        n16880, n16891, n16892, n16595, n16682, n16254, n16253, 
        n16252, n16251, n16250, n555_c, n16819, n16820, n160_adj_1359, 
        n16826, n16832, n454_adj_1361, n16833, n16837, n699_adj_1363, 
        n16838, n650_adj_1366, n16836, n16843, n16844, n506_adj_1370, 
        n16818, n16811, n16594, n16249, n16248, n16247, n166, 
        n16796, n573_c, n16729, n16246, n448_adj_1374, n16862, n16871, 
        n543_c, n16879, n386, n16681, n344_adj_1377, n16890, n16898, 
        n696_adj_1380, n16852, n9531, n16245, n9108, n16244, n16243, 
        n16593, n558_c, n16804, n16805, n16825, n293_adj_1386, n337, 
        n16680;
    wire [14:0]n832_adj_1979;
    
    wire n16831, n16842;
    wire [14:0]n832_adj_1980;
    wire [14:0]n833_adj_1981;
    
    wire n16241, n524, n16728, n16627, n16626, n739_adj_1396, n451_adj_1397, 
        n16847, n16850, n687, n16240, n16861, n16889, n16239, 
        n16238, n16237, n16236, n16235, n16234, n16233, n16232, 
        n16231, n16230, n16229, n16228;
    wire [14:0]n834_adj_1982;
    
    wire n16226, n743_adj_1411, n16225, n16224, n16223, n16222, 
        n16221, n16220, n16219, n16218, n16217, n16216, n16215, 
        n16214, n16213;
    wire [14:0]n835_adj_1983;
    
    wire n16211, n747_adj_1425, n16210, n16209, n16208, n16207, 
        n16206, n16205, n16204, n16203, n16202, n16201, n16200, 
        n16199, n16198;
    wire [14:0]n836_adj_1984;
    
    wire n16196, n751_adj_1446, n16195, n16194, n16193, n16192, 
        n16191, n16190, n16189, n16188, n16187, n16186, n16185, 
        n16184, n16183;
    wire [14:0]n837_adj_1985;
    
    wire n16181, n755_adj_1464, n16180, n16179, n16178, n16177, 
        n16176, n16175, n16174, n16173, n16172, n16171, n16170, 
        n16169, n16168;
    wire [14:0]n838_adj_1986;
    
    wire n16166, n759_adj_1482, n16165, n16164, n16163, n16162, 
        n16161, n16160, n16159, n16158, n16157, n16156, n212_c, 
        n16155, n163, n16154, n16153;
    wire [14:0]n839_adj_1987;
    
    wire n16151, n763_adj_1502, n705, n16150, n656, n16149, n16148, 
        n16147, n509, n16146, n460, n16145, n16144, n362, n16143, 
        n313_adj_1513, n16142, n16141, n215_adj_1517, n16140, n166_adj_1519, 
        n16139, n16138;
    wire [14:0]n840_adj_1988;
    
    wire n16136, n767_adj_1523, n708_adj_1525, n16135, n659_adj_1527, 
        n16134, n16133, n16132, n512_adj_1533, n16131, n463_adj_1535, 
        n16130, n16129, n365_adj_1539, n16128, n316_adj_1541, n16127, 
        n509_adj_1542, n16803, n16126, n218_adj_1546, n16125, n16808, 
        n169_adj_1550, n16124, n16123, n457_adj_1557, n16817;
    wire [14:0]n841_adj_1989;
    
    wire n16121, n771_adj_1561, n711_adj_1563, n16120, n662_adj_1565, 
        n16119, n16118, n16117, n515_adj_1571, n16116, n466_adj_1573, 
        n16115, n16114, n368_adj_1577, n16113, n16835, n16565, n16679, 
        n16564, n16678;
    wire [30:0]n1;
    
    wire n17331, n17330, n17329, n16848, n500_adj_1590, n16849, 
        n157_adj_1592, n16841, n17328, n17327, n17326, n319_adj_1594, 
        n16112, n17325, n17324, n16563, n460_adj_1598, n16802, n705_adj_1600, 
        n16807, n17323, n16816, n356_adj_1605, n16830, n16840, n146_adj_1608, 
        n190, n16677, n16846, n17322, n16111, n17321, n647_adj_1614, 
        n16851, n17320, n16868, n17319, n494_adj_1618, n16878, n17318, 
        n687_adj_1620, n16897, n17317, n17316, n350_adj_1625, n16860, 
        n17315, n16562, n17314, n301_adj_1629, n16859, n17313, n17312, 
        n17311, n17310, n17309, n17308, n17307, n17306, n17305, 
        n97_adj_1633, n16676, n16888, n17304, VCC_net, n221_adj_1638, 
        n16110, n172_adj_1640, n16109, n16108, n16795, n656_adj_1646, 
        n16806, n359_adj_1648, n16815, n638_adj_1649, n16896, n16823, 
        n307_adj_1653, n16829, n552_adj_1654, n16834, n353_adj_1655, 
        n16845, n693_adj_1657, n16867, n16561, n310_adj_1660, n16814, 
        n549_adj_1662, n475, n16727, n16858, n445_adj_1667, n16877, 
        n16876, n48_adj_1670, n16887, n148_adj_1673, n16886, n16560, 
        n16674;
    wire [14:0]n842_adj_1990;
    
    wire n16106, n775_adj_1680, n714_adj_1682, n16105, n665_adj_1684, 
        n16104, n16103, n16102, n518_adj_1690, n16101, n469_adj_1692, 
        n16100, n16099, n371_adj_1696, n16098, n322_adj_1698, n16097, 
        n16096, n224_adj_1702, n16095, n175_adj_1704, n16094, n16093;
    wire [14:0]n843_adj_1991;
    
    wire n16091, n779_adj_1712, n717_adj_1714, n16090, n668_adj_1716, 
        n16089, n16088, n16087, n521_adj_1722, n16086, n472_adj_1724, 
        n16085, n16084, n374_adj_1728, n16083, n325_adj_1730, n16082, 
        n16081, n227_adj_1734, n16080, n178_adj_1736, n16079, n16078;
    wire [14:0]n844_adj_1992;
    
    wire n16076, n783_adj_1744, n720_adj_1746, n16075, n671_adj_1748, 
        n16074, n16073, n347_adj_1751, n16875, n16072, n524_adj_1755, 
        n16071, n475_adj_1757, n16070, n16069, n377, n16068, n328, 
        n16067, n16066, n230_c, n16065, n181, n16064, n16063;
    wire [14:0]n845_adj_1993;
    
    wire n16061, n787_adj_1767, n723_adj_1769, n16060, n674_adj_1771, 
        n16059, n16058, n16057, n16895, n527_adj_1778, n16056, n478_adj_1780, 
        n16055, n16054, n380_adj_1784, n16053, n331_adj_1786, n16052, 
        n16051, n233_adj_1790, n16050, n184_adj_1792, n16049, n16048;
    wire [14:0]n846_adj_1994;
    
    wire n16046, n791_adj_1798, n726, n16045, n677, n16044, n16043, 
        n16042, n530, n16041, n481, n16040, n16039, n383, n16038, 
        n334, n16037, n16036, n236_adj_1810, n16035, n187_adj_1812, 
        n16034, n16033, n19580, n16032, n729_adj_1819, n16031, n636_adj_1820, 
        n680_adj_1821, n16030, n16029, n16028, n533_adj_1827, n16027, 
        n440_adj_1828, n484_adj_1829, n16026, n16025, n386_adj_1833, 
        n16024, n293_adj_1834, n337_adj_1835, n16023, n16022, n239_adj_1839, 
        n16021, n146_adj_1840, n190_adj_1841, n16020, n97_adj_1842, 
        n16019, n48_adj_1844, n16018, n16017, n16016, n16015, n16014, 
        n16013, n16012, n16011, n16010, n16009, n16008, n16007, 
        n16006, n16005, n16004, n17691, n16559, n16673, n16857, 
        n644_adj_1851, n16866, n16885, n377_adj_1853, n17690, n702_adj_1855, 
        n298_adj_1856, n16874, n16558, n16672, n17689, n540_adj_1860, 
        n16894, n16592, n16671, n154_adj_1862, n16813, n16856, n16865, 
        n16873, n16883, n16822, n16557, n16670, n16726, n16725, 
        n16801, n16872, n16893, n151_adj_1886, n690_adj_1887, n442_adj_1889, 
        n653_adj_1891, n16821, n362_adj_1892, n328_adj_1894, n16724, 
        n16812, n17688, n17687, n163_adj_1898, n16548, n16723, n16591, 
        n16669, n16547, n16722, n16549, n181_adj_1904, n16721, n16720, 
        n16590, n16668, n16659, n16667, n16657, n16658, n16666, 
        n16625, n16624, n16665, n16623, n16664, n16718, n723_adj_1912, 
        n16717, n16550, n674_adj_1914, n16716, n17686, n16715, n16551, 
        n576_adj_1918, n16714, n17685, n527_adj_1920, n16713, n17684, 
        n17683, n17682, n17681, n17680, n17679, n17678, n478_adj_1922, 
        n16712, n16711, n16622, n16621, n16620, n16619, n16618, 
        n380_adj_1929, n16710, n331_adj_1931, n16709, n16708, n16707, 
        n184_adj_1935, n16706, n16617, n16616, n16705, n16703, n726_adj_1940, 
        n16702, n677_adj_1941, n16701, n16700, n579_adj_1943, n16699, 
        n530_adj_1944, n16698, n481_adj_1945, n16697, n16696, n383_adj_1947, 
        n16695, n334_adj_1948, n16694, n16663;
    
    SB_LUT4 Q_15__I_0_i210_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n310));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_571_7_lut (.I0(GND_net), .I1(n843[4]), .I2(n331), 
            .I3(n16545), .O(n842[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i369_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n546_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_571_7 (.CI(n16545), .I0(n843[4]), .I1(n331), 
            .CO(n16546));
    SB_LUT4 Q_15__I_0_i243_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n359));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_571_6_lut (.I0(GND_net), .I1(n843[3]), .I2(n282_c), 
            .I3(n16544), .O(n842[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_6 (.CI(n16544), .I0(n843[3]), .I1(n282_c), 
            .CO(n16545));
    SB_LUT4 Q_15__I_0_11_add_571_5_lut (.I0(GND_net), .I1(n843[2]), .I2(n233_c), 
            .I3(n16543), .O(n842[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_5 (.CI(n16543), .I0(n843[2]), .I1(n233_c), 
            .CO(n16544));
    SB_LUT4 Q_15__I_0_11_add_571_4_lut (.I0(GND_net), .I1(n843[1]), .I2(n184), 
            .I3(n16542), .O(n842[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_4 (.CI(n16542), .I0(n843[1]), .I1(n184), 
            .CO(n16543));
    SB_LUT4 Q_15__I_0_11_add_568_5_lut (.I0(GND_net), .I1(n840[2]), .I2(n233_c), 
            .I3(n16588), .O(n839[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_13 (.CI(n16790), .I0(n840_adj_1950[10]), 
            .I1(n610), .CO(n16791));
    SB_CARRY Q_15__I_0_11_add_571_14 (.CI(n16552), .I0(n843[11]), .I1(n674), 
            .CO(n16553));
    SB_LUT4 Q_15__I_0_11_add_571_3_lut (.I0(GND_net), .I1(n843[0]), .I2(n135_c), 
            .I3(n16541), .O(n842[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_i237_2_lut (.I0(\qVoltage[7] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n380));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i309_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i309_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_7655_10 (.CI(n17676), .I0(Product3_mul_temp[10]), .I1(Product4_mul_temp[10]), 
            .CO(n17677));
    SB_CARRY Q_15__I_0_11_add_571_3 (.CI(n16541), .I0(n843[0]), .I1(n135_c), 
            .CO(n16542));
    SB_LUT4 Q_15__I_0_11_add_571_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n842[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16541));
    SB_LUT4 Q_15__I_0_11_add_572_16_lut (.I0(GND_net), .I1(n844[13]), .I2(n793), 
            .I3(n16539), .O(n843[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_16 (.CI(n16539), .I0(n844[13]), .I1(n793), 
            .CO(n783));
    SB_LUT4 Q_15__I_0_11_add_572_15_lut (.I0(GND_net), .I1(n844[12]), .I2(n723), 
            .I3(n16538), .O(n843[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_568_12_lut (.I0(GND_net), .I1(n840_adj_1950[9]), 
            .I2(n561_c), .I3(n16789), .O(n839_adj_1951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_9 (.CI(n17675), .I0(Product3_mul_temp[9]), .I1(Product4_mul_temp[9]), 
            .CO(n17676));
    SB_CARRY Q_15__I_0_11_add_572_15 (.CI(n16538), .I0(n844[12]), .I1(n723), 
            .CO(n16539));
    SB_LUT4 Q_15__I_0_11_add_572_14_lut (.I0(GND_net), .I1(n844[11]), .I2(n674), 
            .I3(n16537), .O(n843[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_8 (.CI(n17674), .I0(Product3_mul_temp[8]), .I1(Product4_mul_temp[8]), 
            .CO(n17675));
    SB_CARRY Q_15__I_0_11_add_572_14 (.CI(n16537), .I0(n844[11]), .I1(n674), 
            .CO(n16538));
    SB_LUT4 Q_15__I_0_11_add_572_13_lut (.I0(GND_net), .I1(n844[10]), .I2(n625_c), 
            .I3(n16536), .O(n843[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_13 (.CI(n16536), .I0(n844[10]), .I1(n625_c), 
            .CO(n16537));
    SB_CARRY D_15__I_0_10_add_568_12 (.CI(n16789), .I0(n840_adj_1950[9]), 
            .I1(n561_c), .CO(n16790));
    SB_LUT4 D_15__I_0_10_i206_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n304));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i342_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n506));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i342_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_572_12_lut (.I0(GND_net), .I1(n844[9]), .I2(n576), 
            .I3(n16535), .O(n843[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_12 (.CI(n16535), .I0(n844[9]), .I1(n576), 
            .CO(n16536));
    SB_LUT4 Q_15__I_0_11_add_572_11_lut (.I0(GND_net), .I1(n844[8]), .I2(n527), 
            .I3(n16534), .O(n843[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_11 (.CI(n16534), .I0(n844[8]), .I1(n527), 
            .CO(n16535));
    SB_CARRY Q_15__I_0_11_add_568_5 (.CI(n16588), .I0(n840[2]), .I1(n233_c), 
            .CO(n16589));
    SB_LUT4 D_15__I_0_10_add_568_11_lut (.I0(GND_net), .I1(n840_adj_1950[8]), 
            .I2(n512), .I3(n16788), .O(n839_adj_1951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_11 (.CI(n16788), .I0(n840_adj_1950[8]), 
            .I1(n512), .CO(n16789));
    SB_LUT4 D_15__I_0_10_add_568_10_lut (.I0(GND_net), .I1(n840_adj_1950[7]), 
            .I2(n463), .I3(n16787), .O(n839_adj_1951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_10 (.CI(n16787), .I0(n840_adj_1950[7]), 
            .I1(n463), .CO(n16788));
    SB_LUT4 D_15__I_0_10_add_568_9_lut (.I0(GND_net), .I1(n840_adj_1950[6]), 
            .I2(n414), .I3(n16786), .O(n839_adj_1951[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_9 (.CI(n16786), .I0(n840_adj_1950[6]), 
            .I1(n414), .CO(n16787));
    SB_LUT4 D_15__I_0_10_add_568_8_lut (.I0(GND_net), .I1(n840_adj_1950[5]), 
            .I2(n365), .I3(n16785), .O(n839_adj_1951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_8 (.CI(n16785), .I0(n840_adj_1950[5]), 
            .I1(n365), .CO(n16786));
    SB_LUT4 D_15__I_0_10_add_568_7_lut (.I0(GND_net), .I1(n840_adj_1950[4]), 
            .I2(n316), .I3(n16784), .O(n839_adj_1951[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_7 (.CI(n16784), .I0(n840_adj_1950[4]), 
            .I1(n316), .CO(n16785));
    SB_LUT4 D_15__I_0_10_add_568_6_lut (.I0(GND_net), .I1(n840_adj_1950[3]), 
            .I2(n267), .I3(n16783), .O(n839_adj_1951[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_6 (.CI(n16783), .I0(n840_adj_1950[3]), 
            .I1(n267), .CO(n16784));
    SB_LUT4 D_15__I_0_10_add_568_5_lut (.I0(GND_net), .I1(n840_adj_1950[2]), 
            .I2(n218), .I3(n16782), .O(n839_adj_1951[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_5 (.CI(n16782), .I0(n840_adj_1950[2]), 
            .I1(n218), .CO(n16783));
    SB_CARRY Q_15__I_0_11_add_564_12 (.CI(n16655), .I0(n836[9]), .I1(n576), 
            .CO(n16656));
    SB_LUT4 Q_15__I_0_i441_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n653));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i441_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i474_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n702));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i474_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i402_2_lut (.I0(\qVoltage[12] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n625_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_574_5 (.CI(n16692), .I0(n846[2]), .I1(n236), 
            .CO(n16693));
    SB_LUT4 D_15__I_0_10_add_568_4_lut (.I0(GND_net), .I1(n840_adj_1950[1]), 
            .I2(n169), .I3(n16781), .O(n839_adj_1951[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_568_4_lut (.I0(GND_net), .I1(n840[1]), .I2(n184), 
            .I3(n16587), .O(n839[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_11_lut (.I0(GND_net), .I1(n836[8]), .I2(n527), 
            .I3(n16654), .O(n835[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_4 (.CI(n16781), .I0(n840_adj_1950[1]), 
            .I1(n169), .CO(n16782));
    SB_CARRY add_7655_7 (.CI(n17673), .I0(Product3_mul_temp[7]), .I1(Product4_mul_temp[7]), 
            .CO(n17674));
    SB_CARRY Q_15__I_0_11_add_564_11 (.CI(n16654), .I0(n836[8]), .I1(n527), 
            .CO(n16655));
    SB_LUT4 D_15__I_0_10_add_568_3_lut (.I0(GND_net), .I1(n840_adj_1950[0]), 
            .I2(n120), .I3(n16780), .O(n839_adj_1951[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i109_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n160));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_564_10_lut (.I0(GND_net), .I1(n836[7]), .I2(n478), 
            .I3(n16653), .O(n835[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i332_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n491));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i332_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_7655_6 (.CI(n17672), .I0(Product3_mul_temp[6]), .I1(Product4_mul_temp[6]), 
            .CO(n17673));
    SB_LUT4 Q_15__I_0_i142_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n209_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i208_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n307));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i241_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n356));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i241_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_568_3 (.CI(n16780), .I0(n840_adj_1950[0]), 
            .I1(n120), .CO(n16781));
    SB_CARRY add_7655_5 (.CI(n17671), .I0(Product3_mul_temp[5]), .I1(Product4_mul_temp[5]), 
            .CO(n17672));
    SB_CARRY add_7655_4 (.CI(n17670), .I0(Product3_mul_temp[4]), .I1(Product4_mul_temp[4]), 
            .CO(n17671));
    SB_CARRY add_7655_3 (.CI(n17669), .I0(Product3_mul_temp[3]), .I1(Product4_mul_temp[3]), 
            .CO(n17670));
    SB_CARRY add_7655_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), .I1(Product4_mul_temp[2]), 
            .CO(n17669));
    SB_LUT4 Q_15__I_0_11_add_572_10_lut (.I0(GND_net), .I1(n844[7]), .I2(n478), 
            .I3(n16533), .O(n843[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_568_2_lut (.I0(GND_net), .I1(n26), .I2(n71), 
            .I3(GND_net), .O(n839_adj_1951[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_574_4_lut (.I0(GND_net), .I1(n846[1]), .I2(n187), 
            .I3(n16691), .O(n845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_3_lut (.I0(GND_net), .I1(n835[0]), .I2(n135_c), 
            .I3(n16661), .O(Product2_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_4 (.CI(n16691), .I0(n846[1]), .I1(n187), 
            .CO(n16692));
    SB_CARRY Q_15__I_0_11_add_570_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16556));
    SB_LUT4 D_15__I_0_10_add_574_3_lut (.I0(GND_net), .I1(n846[0]), .I2(n138), 
            .I3(n16690), .O(n845[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_3 (.CI(n16661), .I0(n835[0]), .I1(n135_c), 
            .CO(n16662));
    SB_CARRY D_15__I_0_10_add_574_3 (.CI(n16690), .I0(n846[0]), .I1(n138), 
            .CO(n16691));
    SB_LUT4 D_15__I_0_10_add_574_2_lut (.I0(GND_net), .I1(n44), .I2(n89), 
            .I3(GND_net), .O(n845[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16661));
    SB_LUT4 add_7655_30_lut (.I0(GND_net), .I1(Product3_mul_temp[29]), .I2(Product4_mul_temp[29]), 
            .I3(n17696), .O(\betaVoltage[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_5 (.CI(n16827), .I0(n837[2]), .I1(n209), 
            .CO(n16828));
    SB_CARRY Q_15__I_0_11_add_572_10 (.CI(n16533), .I0(n844[7]), .I1(n478), 
            .CO(n16534));
    SB_CARRY D_15__I_0_10_add_574_2 (.CI(GND_net), .I0(n44), .I1(n89), 
            .CO(n16690));
    SB_CARRY D_15__I_0_10_add_568_2 (.CI(GND_net), .I0(n26), .I1(n71), 
            .CO(n16780));
    SB_CARRY Q_15__I_0_11_add_564_10 (.CI(n16653), .I0(n836[7]), .I1(n478), 
            .CO(n16654));
    SB_LUT4 Q_15__I_0_11_add_568_3_lut (.I0(GND_net), .I1(n840[0]), .I2(n135_c), 
            .I3(n16586), .O(n839[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_568_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n839[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7655_29_lut (.I0(GND_net), .I1(Product3_mul_temp[29]), .I2(Product4_mul_temp[29]), 
            .I3(n17695), .O(\betaVoltage[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_16_lut (.I0(GND_net), .I1(n19681), .I2(n19684), 
            .I3(n16689), .O(n846[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_3 (.CI(n16586), .I0(n840[0]), .I1(n135_c), 
            .CO(n16587));
    SB_LUT4 D_15__I_0_10_add_569_16_lut (.I0(GND_net), .I1(n841[13]), .I2(n769), 
            .I3(n16778), .O(n840_adj_1950[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_16 (.CI(n16554), .I0(n843[13]), .I1(n793), 
            .CO(n779));
    SB_LUT4 Q_15__I_0_11_add_572_9_lut (.I0(GND_net), .I1(n844[6]), .I2(n429_c), 
            .I3(n16532), .O(n843[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i307_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i307_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_572_9 (.CI(n16532), .I0(n844[6]), .I1(n429_c), 
            .CO(n16533));
    SB_LUT4 Q_15__I_0_11_add_572_8_lut (.I0(GND_net), .I1(n844[5]), .I2(n380), 
            .I3(n16531), .O(n843[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i340_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n503));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i340_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_569_16 (.CI(n16778), .I0(n841[13]), .I1(n769), 
            .CO(n771));
    SB_CARRY add_7655_29 (.CI(n17695), .I0(Product3_mul_temp[29]), .I1(Product4_mul_temp[29]), 
            .CO(n17696));
    SB_CARRY Q_15__I_0_11_add_568_4 (.CI(n16587), .I0(n840[1]), .I1(n184), 
            .CO(n16588));
    SB_LUT4 D_15__I_0_10_add_575_15_lut (.I0(GND_net), .I1(n685), .I2(n729), 
            .I3(n16688), .O(n846[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16586));
    SB_CARRY D_15__I_0_10_add_575_15 (.CI(n16688), .I0(n685), .I1(n729), 
            .CO(n16689));
    SB_LUT4 Q_15__I_0_11_add_569_16_lut (.I0(GND_net), .I1(n841_adj_1952[13]), 
            .I2(n793), .I3(n16584), .O(n840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_14_lut (.I0(GND_net), .I1(n636), .I2(n680), 
            .I3(n16687), .O(n846[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_16 (.CI(n16584), .I0(n841_adj_1952[13]), 
            .I1(n793), .CO(n771_adj_1019));
    SB_CARRY D_15__I_0_10_add_575_14 (.CI(n16687), .I0(n636), .I1(n680), 
            .CO(n16688));
    SB_LUT4 D_15__I_0_10_add_569_15_lut (.I0(GND_net), .I1(n841[12]), .I2(n711), 
            .I3(n16777), .O(n840_adj_1950[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_15 (.CI(n16777), .I0(n841[12]), .I1(n711), 
            .CO(n16778));
    SB_LUT4 D_15__I_0_10_add_575_13_lut (.I0(GND_net), .I1(n587), .I2(n631), 
            .I3(n16686), .O(n846[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_569_14_lut (.I0(GND_net), .I1(n841[11]), .I2(n662), 
            .I3(n16776), .O(n840_adj_1950[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7655_28_lut (.I0(GND_net), .I1(Product3_mul_temp[28]), .I2(Product4_mul_temp[28]), 
            .I3(n17694), .O(\betaVoltage[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i340_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n503_adj_1020));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i340_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_567_7 (.CI(n16799), .I0(n839_adj_1951[4]), 
            .I1(n313), .CO(n16800));
    SB_CARRY Q_15__I_0_11_add_572_8 (.CI(n16531), .I0(n844[5]), .I1(n380), 
            .CO(n16532));
    SB_LUT4 D_15__I_0_10_add_567_6_lut (.I0(GND_net), .I1(n839_adj_1951[3]), 
            .I2(n264), .I3(n16798), .O(n838[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_566_3_lut (.I0(GND_net), .I1(n838[0]), .I2(n114), 
            .I3(n16810), .O(n837[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_15 (.CI(n16792), .I0(n840_adj_1950[12]), 
            .I1(n708), .CO(n16793));
    SB_LUT4 Q_15__I_0_11_add_572_7_lut (.I0(GND_net), .I1(n844[4]), .I2(n331), 
            .I3(n16530), .O(n843[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_14 (.CI(n16776), .I0(n841[11]), .I1(n662), 
            .CO(n16777));
    SB_CARRY Q_15__I_0_11_add_569_15 (.CI(n16583), .I0(n841_adj_1952[12]), 
            .I1(n723), .CO(n16584));
    SB_LUT4 Q_15__I_0_11_add_569_15_lut (.I0(GND_net), .I1(n841_adj_1952[12]), 
            .I2(n723), .I3(n16583), .O(n840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i439_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n650));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i439_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_567_14_lut (.I0(GND_net), .I1(n839[11]), .I2(n674), 
            .I3(n16612), .O(n838_adj_1953[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_15 (.CI(n16613), .I0(n839[12]), .I1(n723), 
            .CO(n16614));
    SB_LUT4 Q_15__I_0_i472_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n699));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i472_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_567_13 (.CI(n16611), .I0(n839[10]), .I1(n625_c), 
            .CO(n16612));
    SB_LUT4 Q_15__I_0_11_add_567_13_lut (.I0(GND_net), .I1(n839[10]), .I2(n625_c), 
            .I3(n16611), .O(n838_adj_1953[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_14 (.CI(n16612), .I0(n839[11]), .I1(n674), 
            .CO(n16613));
    SB_LUT4 Q_15__I_0_11_add_569_14_lut (.I0(GND_net), .I1(n841_adj_1952[11]), 
            .I2(n674), .I3(n16582), .O(n840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_567_12_lut (.I0(GND_net), .I1(n839[9]), .I2(n576), 
            .I3(n16610), .O(n838_adj_1953[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_12 (.CI(n16610), .I0(n839[9]), .I1(n576), 
            .CO(n16611));
    SB_CARRY Q_15__I_0_11_add_567_11 (.CI(n16609), .I0(n839[8]), .I1(n527), 
            .CO(n16610));
    SB_LUT4 Q_15__I_0_11_add_567_11_lut (.I0(GND_net), .I1(n839[8]), .I2(n527), 
            .I3(n16609), .O(n838_adj_1953[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_567_10_lut (.I0(GND_net), .I1(n839[7]), .I2(n478), 
            .I3(n16608), .O(n838_adj_1953[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_9_lut (.I0(GND_net), .I1(n836[6]), .I2(n429_c), 
            .I3(n16652), .O(n835[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_569_13_lut (.I0(GND_net), .I1(n841[10]), .I2(n613), 
            .I3(n16775), .O(n840_adj_1950[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_13 (.CI(n16775), .I0(n841[10]), .I1(n613), 
            .CO(n16776));
    SB_LUT4 D_15__I_0_10_add_569_12_lut (.I0(GND_net), .I1(n841[9]), .I2(n564_c), 
            .I3(n16774), .O(n840_adj_1950[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i107_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n157));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i107_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_564_9 (.CI(n16652), .I0(n836[6]), .I1(n429_c), 
            .CO(n16653));
    SB_CARRY D_15__I_0_10_add_569_12 (.CI(n16774), .I0(n841[9]), .I1(n564_c), 
            .CO(n16775));
    SB_LUT4 D_15__I_0_10_add_569_11_lut (.I0(GND_net), .I1(n841[8]), .I2(n515), 
            .I3(n16773), .O(n840_adj_1950[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i379_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n561_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_564_8_lut (.I0(GND_net), .I1(n836[5]), .I2(n380), 
            .I3(n16651), .O(n835[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_11 (.CI(n16773), .I0(n841[8]), .I1(n515), 
            .CO(n16774));
    SB_LUT4 D_15__I_0_10_add_569_10_lut (.I0(GND_net), .I1(n841[7]), .I2(n466), 
            .I3(n16772), .O(n840_adj_1950[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_10 (.CI(n16772), .I0(n841[7]), .I1(n466), 
            .CO(n16773));
    SB_CARRY Q_15__I_0_11_add_564_8 (.CI(n16651), .I0(n836[5]), .I1(n380), 
            .CO(n16652));
    SB_LUT4 D_15__I_0_10_add_569_9_lut (.I0(GND_net), .I1(n841[6]), .I2(n417), 
            .I3(n16771), .O(n840_adj_1950[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_7_lut (.I0(GND_net), .I1(n836[4]), .I2(n331), 
            .I3(n16650), .O(n835[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_9 (.CI(n16771), .I0(n841[6]), .I1(n417), 
            .CO(n16772));
    SB_CARRY Q_15__I_0_11_add_564_7 (.CI(n16650), .I0(n836[4]), .I1(n331), 
            .CO(n16651));
    SB_LUT4 Q_15__I_0_i140_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n206_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_add_569_8_lut (.I0(GND_net), .I1(n841[5]), .I2(n368), 
            .I3(n16770), .O(n840_adj_1950[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_6_lut (.I0(GND_net), .I1(n836[3]), .I2(n282_c), 
            .I3(n16649), .O(n835[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_8 (.CI(n16770), .I0(n841[5]), .I1(n368), 
            .CO(n16771));
    SB_LUT4 D_15__I_0_10_add_569_7_lut (.I0(GND_net), .I1(n841[4]), .I2(n319), 
            .I3(n16769), .O(n840_adj_1950[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_564_6 (.CI(n16649), .I0(n836[3]), .I1(n282_c), 
            .CO(n16650));
    SB_CARRY D_15__I_0_10_add_569_7 (.CI(n16769), .I0(n841[4]), .I1(n319), 
            .CO(n16770));
    SB_CARRY add_7655_28 (.CI(n17694), .I0(Product3_mul_temp[28]), .I1(Product4_mul_temp[28]), 
            .CO(n17695));
    SB_LUT4 Q_15__I_0_11_add_569_13_lut (.I0(GND_net), .I1(n841_adj_1952[10]), 
            .I2(n625_c), .I3(n16581), .O(n840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_14 (.CI(n16582), .I0(n841_adj_1952[11]), 
            .I1(n674), .CO(n16583));
    SB_LUT4 Q_15__I_0_i206_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n304_adj_1031));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_567_9_lut (.I0(GND_net), .I1(n839[6]), .I2(n429_c), 
            .I3(n16607), .O(n838_adj_1953[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_10 (.CI(n16608), .I0(n839[7]), .I1(n478), 
            .CO(n16609));
    SB_CARRY Q_15__I_0_11_add_567_8 (.CI(n16606), .I0(n839[5]), .I1(n380), 
            .CO(n16607));
    SB_LUT4 Q_15__I_0_11_add_567_8_lut (.I0(GND_net), .I1(n839[5]), .I2(n380), 
            .I3(n16606), .O(n838_adj_1953[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_9 (.CI(n16607), .I0(n839[6]), .I1(n429_c), 
            .CO(n16608));
    SB_CARRY Q_15__I_0_11_add_569_13 (.CI(n16581), .I0(n841_adj_1952[10]), 
            .I1(n625_c), .CO(n16582));
    SB_LUT4 Q_15__I_0_i239_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n353));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_567_7_lut (.I0(GND_net), .I1(n839[4]), .I2(n331), 
            .I3(n16605), .O(n838_adj_1953[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i305_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i305_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_567_7 (.CI(n16605), .I0(n839[4]), .I1(n331), 
            .CO(n16606));
    SB_LUT4 add_7655_27_lut (.I0(GND_net), .I1(Product3_mul_temp[27]), .I2(Product4_mul_temp[27]), 
            .I3(n17693), .O(\betaVoltage[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i338_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n500));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i338_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_567_6 (.CI(n16604), .I0(n839[3]), .I1(n282_c), 
            .CO(n16605));
    SB_LUT4 Q_15__I_0_11_add_567_6_lut (.I0(GND_net), .I1(n839[3]), .I2(n282_c), 
            .I3(n16604), .O(n838_adj_1953[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_567_5_lut (.I0(GND_net), .I1(n839[2]), .I2(n233_c), 
            .I3(n16603), .O(n838_adj_1953[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_i270_2_lut (.I0(\qVoltage[8] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n429_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_564_5_lut (.I0(GND_net), .I1(n836[2]), .I2(n233_c), 
            .I3(n16648), .O(n835[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_569_6_lut (.I0(GND_net), .I1(n841[3]), .I2(n270), 
            .I3(n16768), .O(n840_adj_1950[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_6 (.CI(n16768), .I0(n841[3]), .I1(n270), 
            .CO(n16769));
    SB_LUT4 D_15__I_0_10_add_569_5_lut (.I0(GND_net), .I1(n841[2]), .I2(n221), 
            .I3(n16767), .O(n840_adj_1950[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_564_5 (.CI(n16648), .I0(n836[2]), .I1(n233_c), 
            .CO(n16649));
    SB_CARRY D_15__I_0_10_add_569_5 (.CI(n16767), .I0(n841[2]), .I1(n221), 
            .CO(n16768));
    SB_LUT4 D_15__I_0_10_add_569_4_lut (.I0(GND_net), .I1(n841[1]), .I2(n172), 
            .I3(n16766), .O(n840_adj_1950[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_4_lut (.I0(GND_net), .I1(n836[1]), .I2(n184), 
            .I3(n16647), .O(n835[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_4 (.CI(n16766), .I0(n841[1]), .I1(n172), 
            .CO(n16767));
    SB_LUT4 D_15__I_0_10_add_569_3_lut (.I0(GND_net), .I1(n841[0]), .I2(n123), 
            .I3(n16765), .O(n840_adj_1950[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_3 (.CI(n16765), .I0(n841[0]), .I1(n123), 
            .CO(n16766));
    SB_CARRY Q_15__I_0_11_add_564_4 (.CI(n16647), .I0(n836[1]), .I1(n184), 
            .CO(n16648));
    SB_LUT4 D_15__I_0_10_add_569_2_lut (.I0(GND_net), .I1(n29), .I2(n74), 
            .I3(GND_net), .O(n840_adj_1950[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_3_lut (.I0(GND_net), .I1(n836[0]), .I2(n135_c), 
            .I3(n16646), .O(n835[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_569_2 (.CI(GND_net), .I0(n29), .I1(n74), 
            .CO(n16765));
    SB_LUT4 Q_15__I_0_i437_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n647));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i437_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i470_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n696));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i470_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_564_3 (.CI(n16646), .I0(n836[0]), .I1(n135_c), 
            .CO(n16647));
    SB_LUT4 D_15__I_0_10_add_570_16_lut (.I0(GND_net), .I1(n842_adj_1954[13]), 
            .I2(n773), .I3(n16763), .O(n841[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n835[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_16 (.CI(n16763), .I0(n842_adj_1954[13]), 
            .I1(n773), .CO(n775));
    SB_LUT4 D_15__I_0_10_add_570_15_lut (.I0(GND_net), .I1(n842_adj_1954[12]), 
            .I2(n714), .I3(n16762), .O(n841[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_564_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16646));
    SB_CARRY D_15__I_0_10_add_570_15 (.CI(n16762), .I0(n842_adj_1954[12]), 
            .I1(n714), .CO(n16763));
    SB_CARRY Q_15__I_0_11_add_572_7 (.CI(n16530), .I0(n844[4]), .I1(n331), 
            .CO(n16531));
    SB_LUT4 Q_15__I_0_11_add_565_16_lut (.I0(GND_net), .I1(n837_adj_1955[13]), 
            .I2(n793), .I3(n16644), .O(n836[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_570_14_lut (.I0(GND_net), .I1(n842_adj_1954[11]), 
            .I2(n665), .I3(n16761), .O(n841[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_14 (.CI(n16761), .I0(n842_adj_1954[11]), 
            .I1(n665), .CO(n16762));
    SB_LUT4 D_15__I_0_10_add_570_13_lut (.I0(GND_net), .I1(n842_adj_1954[10]), 
            .I2(n616), .I3(n16760), .O(n841[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_13 (.CI(n16760), .I0(n842_adj_1954[10]), 
            .I1(n616), .CO(n16761));
    SB_LUT4 D_15__I_0_10_add_570_12_lut (.I0(GND_net), .I1(n842_adj_1954[9]), 
            .I2(n567_c), .I3(n16759), .O(n841[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_12 (.CI(n16759), .I0(n842_adj_1954[9]), 
            .I1(n567_c), .CO(n16760));
    SB_LUT4 D_15__I_0_10_add_570_11_lut (.I0(GND_net), .I1(n842_adj_1954[8]), 
            .I2(n518), .I3(n16758), .O(n841[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_11 (.CI(n16758), .I0(n842_adj_1954[8]), 
            .I1(n518), .CO(n16759));
    SB_LUT4 D_15__I_0_10_add_570_10_lut (.I0(GND_net), .I1(n842_adj_1954[7]), 
            .I2(n469), .I3(n16757), .O(n841[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_10 (.CI(n16757), .I0(n842_adj_1954[7]), 
            .I1(n469), .CO(n16758));
    SB_LUT4 D_15__I_0_10_add_570_9_lut (.I0(GND_net), .I1(n842_adj_1954[6]), 
            .I2(n420), .I3(n16756), .O(n841[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_9 (.CI(n16756), .I0(n842_adj_1954[6]), 
            .I1(n420), .CO(n16757));
    SB_LUT4 Q_15__I_0_i105_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n154));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i105_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_7655_27 (.CI(n17693), .I0(Product3_mul_temp[27]), .I1(Product4_mul_temp[27]), 
            .CO(n17694));
    SB_CARRY Q_15__I_0_11_add_569_9 (.CI(n16577), .I0(n841_adj_1952[6]), 
            .I1(n429_c), .CO(n16578));
    SB_LUT4 Q_15__I_0_11_add_569_9_lut (.I0(GND_net), .I1(n841_adj_1952[6]), 
            .I2(n429_c), .I3(n16577), .O(n840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_10 (.CI(n16578), .I0(n841_adj_1952[7]), 
            .I1(n478), .CO(n16579));
    SB_LUT4 Q_15__I_0_11_add_569_10_lut (.I0(GND_net), .I1(n841_adj_1952[7]), 
            .I2(n478), .I3(n16578), .O(n840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_11 (.CI(n16579), .I0(n841_adj_1952[8]), 
            .I1(n527), .CO(n16580));
    SB_LUT4 Q_15__I_0_11_add_569_11_lut (.I0(GND_net), .I1(n841_adj_1952[8]), 
            .I2(n527), .I3(n16579), .O(n840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_12 (.CI(n16580), .I0(n841_adj_1952[9]), 
            .I1(n576), .CO(n16581));
    SB_LUT4 Q_15__I_0_11_add_569_12_lut (.I0(GND_net), .I1(n841_adj_1952[9]), 
            .I2(n576), .I3(n16580), .O(n840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i138_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n203_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i138_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_567_5 (.CI(n16603), .I0(n839[2]), .I1(n233_c), 
            .CO(n16604));
    SB_LUT4 Q_15__I_0_11_add_567_4_lut (.I0(GND_net), .I1(n839[1]), .I2(n184), 
            .I3(n16602), .O(n838_adj_1953[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7655_26_lut (.I0(GND_net), .I1(Product3_mul_temp[26]), .I2(Product4_mul_temp[26]), 
            .I3(n17692), .O(\betaVoltage[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_567_3_lut (.I0(GND_net), .I1(n839[0]), .I2(n135_c), 
            .I3(n16601), .O(n838_adj_1953[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_4 (.CI(n16602), .I0(n839[1]), .I1(n184), 
            .CO(n16603));
    SB_CARRY Q_15__I_0_11_add_567_3 (.CI(n16601), .I0(n839[0]), .I1(n135_c), 
            .CO(n16602));
    SB_LUT4 Q_15__I_0_i204_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n301));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i237_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n350));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i237_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_569_6 (.CI(n16574), .I0(n841_adj_1952[3]), 
            .I1(n282_c), .CO(n16575));
    SB_LUT4 Q_15__I_0_11_add_569_6_lut (.I0(GND_net), .I1(n841_adj_1952[3]), 
            .I2(n282_c), .I3(n16574), .O(n840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_7 (.CI(n16575), .I0(n841_adj_1952[4]), 
            .I1(n331), .CO(n16576));
    SB_LUT4 Q_15__I_0_11_add_569_7_lut (.I0(GND_net), .I1(n841_adj_1952[4]), 
            .I2(n331), .I3(n16575), .O(n840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_8 (.CI(n16576), .I0(n841_adj_1952[5]), 
            .I1(n380), .CO(n16577));
    SB_LUT4 Q_15__I_0_11_add_569_8_lut (.I0(GND_net), .I1(n841_adj_1952[5]), 
            .I2(n380), .I3(n16576), .O(n840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i303_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i303_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i336_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n497));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i336_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_565_16 (.CI(n16644), .I0(n837_adj_1955[13]), 
            .I1(n793), .CO(n755));
    SB_LUT4 D_15__I_0_10_add_570_8_lut (.I0(GND_net), .I1(n842_adj_1954[5]), 
            .I2(n371), .I3(n16755), .O(n841[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_15_lut (.I0(GND_net), .I1(n837_adj_1955[12]), 
            .I2(n723), .I3(n16643), .O(n836[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_8 (.CI(n16755), .I0(n842_adj_1954[5]), 
            .I1(n371), .CO(n16756));
    SB_CARRY Q_15__I_0_11_add_565_15 (.CI(n16643), .I0(n837_adj_1955[12]), 
            .I1(n723), .CO(n16644));
    SB_LUT4 D_15__I_0_10_add_570_7_lut (.I0(GND_net), .I1(n842_adj_1954[4]), 
            .I2(n322), .I3(n16754), .O(n841[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_7 (.CI(n16754), .I0(n842_adj_1954[4]), 
            .I1(n322), .CO(n16755));
    SB_LUT4 Q_15__I_0_11_add_565_14_lut (.I0(GND_net), .I1(n837_adj_1955[11]), 
            .I2(n674), .I3(n16642), .O(n836[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_570_6_lut (.I0(GND_net), .I1(n842_adj_1954[3]), 
            .I2(n273), .I3(n16753), .O(n841[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_14 (.CI(n16642), .I0(n837_adj_1955[11]), 
            .I1(n674), .CO(n16643));
    SB_CARRY D_15__I_0_10_add_570_6 (.CI(n16753), .I0(n842_adj_1954[3]), 
            .I1(n273), .CO(n16754));
    SB_LUT4 D_15__I_0_10_add_570_5_lut (.I0(GND_net), .I1(n842_adj_1954[2]), 
            .I2(n224), .I3(n16752), .O(n841[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_5 (.CI(n16752), .I0(n842_adj_1954[2]), 
            .I1(n224), .CO(n16753));
    SB_LUT4 D_15__I_0_10_add_570_4_lut (.I0(GND_net), .I1(n842_adj_1954[1]), 
            .I2(n175), .I3(n16751), .O(n841[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_4 (.CI(n16751), .I0(n842_adj_1954[1]), 
            .I1(n175), .CO(n16752));
    SB_LUT4 D_15__I_0_10_add_570_3_lut (.I0(GND_net), .I1(n842_adj_1954[0]), 
            .I2(n126), .I3(n16750), .O(n841[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16571));
    SB_LUT4 Q_15__I_0_11_add_569_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_3 (.CI(n16571), .I0(n841_adj_1952[0]), 
            .I1(n135_c), .CO(n16572));
    SB_LUT4 Q_15__I_0_11_add_569_3_lut (.I0(GND_net), .I1(n841_adj_1952[0]), 
            .I2(n135_c), .I3(n16571), .O(n840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_4 (.CI(n16572), .I0(n841_adj_1952[1]), 
            .I1(n184), .CO(n16573));
    SB_LUT4 Q_15__I_0_11_add_569_4_lut (.I0(GND_net), .I1(n841_adj_1952[1]), 
            .I2(n184), .I3(n16572), .O(n840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_569_5 (.CI(n16573), .I0(n841_adj_1952[2]), 
            .I1(n233_c), .CO(n16574));
    SB_LUT4 Q_15__I_0_11_add_569_5_lut (.I0(GND_net), .I1(n841_adj_1952[2]), 
            .I2(n233_c), .I3(n16573), .O(n840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_26 (.CI(n17692), .I0(Product3_mul_temp[26]), .I1(Product4_mul_temp[26]), 
            .CO(n17693));
    SB_LUT4 Q_15__I_0_11_add_567_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n838_adj_1953[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16601));
    SB_LUT4 Q_15__I_0_i435_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n644));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i435_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_568_16 (.CI(n16599), .I0(n840[13]), .I1(n793), 
            .CO(n767));
    SB_LUT4 Q_15__I_0_11_add_568_16_lut (.I0(GND_net), .I1(n840[13]), .I2(n793), 
            .I3(n16599), .O(n839[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i468_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n693));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_568_15_lut (.I0(GND_net), .I1(n840[12]), .I2(n723), 
            .I3(n16598), .O(n839[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_14 (.CI(n16567), .I0(n842[11]), .I1(n674), 
            .CO(n16568));
    SB_LUT4 Q_15__I_0_11_add_570_14_lut (.I0(GND_net), .I1(n842[11]), .I2(n674), 
            .I3(n16567), .O(n841_adj_1952[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_15 (.CI(n16568), .I0(n842[12]), .I1(n723), 
            .CO(n16569));
    SB_LUT4 Q_15__I_0_11_add_570_15_lut (.I0(GND_net), .I1(n842[12]), .I2(n723), 
            .I3(n16568), .O(n841_adj_1952[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_16 (.CI(n16569), .I0(n842[13]), .I1(n793), 
            .CO(n775_adj_1064));
    SB_LUT4 Q_15__I_0_11_add_570_16_lut (.I0(GND_net), .I1(n842[13]), .I2(n793), 
            .I3(n16569), .O(n841_adj_1952[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_13_lut (.I0(GND_net), .I1(n837_adj_1955[10]), 
            .I2(n625_c), .I3(n16641), .O(n836[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_3 (.CI(n16750), .I0(n842_adj_1954[0]), 
            .I1(n126), .CO(n16751));
    SB_CARRY Q_15__I_0_11_add_565_13 (.CI(n16641), .I0(n837_adj_1955[10]), 
            .I1(n625_c), .CO(n16642));
    SB_LUT4 D_15__I_0_10_add_570_2_lut (.I0(GND_net), .I1(n32), .I2(n77), 
            .I3(GND_net), .O(n841[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_12_lut (.I0(GND_net), .I1(n837_adj_1955[9]), 
            .I2(n576), .I3(n16640), .O(n836[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_570_2 (.CI(GND_net), .I0(n32), .I1(n77), 
            .CO(n16750));
    SB_LUT4 D_15__I_0_10_add_571_16_lut (.I0(GND_net), .I1(n843_adj_1956[13]), 
            .I2(n777), .I3(n16748), .O(n842_adj_1954[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_12 (.CI(n16640), .I0(n837_adj_1955[9]), 
            .I1(n576), .CO(n16641));
    SB_CARRY D_15__I_0_10_add_571_16 (.CI(n16748), .I0(n843_adj_1956[13]), 
            .I1(n777), .CO(n779_adj_1067));
    SB_LUT4 Q_15__I_0_11_add_565_11_lut (.I0(GND_net), .I1(n837_adj_1955[8]), 
            .I2(n527), .I3(n16639), .O(n836[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_15_lut (.I0(GND_net), .I1(n843_adj_1956[12]), 
            .I2(n717), .I3(n16747), .O(n842_adj_1954[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_15 (.CI(n16747), .I0(n843_adj_1956[12]), 
            .I1(n717), .CO(n16748));
    SB_LUT4 D_15__I_0_10_add_571_14_lut (.I0(GND_net), .I1(n843_adj_1956[11]), 
            .I2(n668), .I3(n16746), .O(n842_adj_1954[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_14 (.CI(n16746), .I0(n843_adj_1956[11]), 
            .I1(n668), .CO(n16747));
    SB_LUT4 D_15__I_0_10_add_571_13_lut (.I0(GND_net), .I1(n843_adj_1956[10]), 
            .I2(n619), .I3(n16745), .O(n842_adj_1954[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_13 (.CI(n16745), .I0(n843_adj_1956[10]), 
            .I1(n619), .CO(n16746));
    SB_LUT4 Q_15__I_0_11_add_572_6_lut (.I0(GND_net), .I1(n844[3]), .I2(n282_c), 
            .I3(n16529), .O(n843[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_6 (.CI(n16529), .I0(n844[3]), .I1(n282_c), 
            .CO(n16530));
    SB_CARRY Q_15__I_0_11_add_565_11 (.CI(n16639), .I0(n837_adj_1955[8]), 
            .I1(n527), .CO(n16640));
    SB_LUT4 Q_15__I_0_11_add_572_5_lut (.I0(GND_net), .I1(n844[2]), .I2(n233_c), 
            .I3(n16528), .O(n843[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_12_lut (.I0(GND_net), .I1(n843_adj_1956[9]), 
            .I2(n570_c), .I3(n16744), .O(n842_adj_1954[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_10_lut (.I0(GND_net), .I1(n837_adj_1955[7]), 
            .I2(n478), .I3(n16638), .O(n836[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_10 (.CI(n16638), .I0(n837_adj_1955[7]), 
            .I1(n478), .CO(n16639));
    SB_LUT4 Q_15__I_0_11_add_565_9_lut (.I0(GND_net), .I1(n837_adj_1955[6]), 
            .I2(n429_c), .I3(n16637), .O(n836[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_5 (.CI(n16528), .I0(n844[2]), .I1(n233_c), 
            .CO(n16529));
    SB_LUT4 Q_15__I_0_11_add_572_4_lut (.I0(GND_net), .I1(n844[1]), .I2(n184), 
            .I3(n16527), .O(n843[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_4 (.CI(n16527), .I0(n844[1]), .I1(n184), 
            .CO(n16528));
    SB_LUT4 Q_15__I_0_11_add_572_3_lut (.I0(GND_net), .I1(n844[0]), .I2(n135_c), 
            .I3(n16526), .O(n843[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_3 (.CI(n16526), .I0(n844[0]), .I1(n135_c), 
            .CO(n16527));
    SB_LUT4 Q_15__I_0_11_add_572_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n843[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_572_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16526));
    SB_LUT4 Q_15__I_0_11_add_573_16_lut (.I0(GND_net), .I1(n845_adj_1957[13]), 
            .I2(n793), .I3(n16524), .O(n844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_16 (.CI(n16524), .I0(n845_adj_1957[13]), 
            .I1(n793), .CO(n787));
    SB_LUT4 Q_15__I_0_11_add_573_15_lut (.I0(GND_net), .I1(n845_adj_1957[12]), 
            .I2(n723), .I3(n16523), .O(n844[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_15 (.CI(n16523), .I0(n845_adj_1957[12]), 
            .I1(n723), .CO(n16524));
    SB_LUT4 Q_15__I_0_11_add_573_14_lut (.I0(GND_net), .I1(n845_adj_1957[11]), 
            .I2(n674), .I3(n16522), .O(n844[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i103_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n151));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i103_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_573_14 (.CI(n16522), .I0(n845_adj_1957[11]), 
            .I1(n674), .CO(n16523));
    SB_LUT4 Q_15__I_0_11_add_573_13_lut (.I0(GND_net), .I1(n845_adj_1957[10]), 
            .I2(n625_c), .I3(n16521), .O(n844[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_13 (.CI(n16521), .I0(n845_adj_1957[10]), 
            .I1(n625_c), .CO(n16522));
    SB_LUT4 Q_15__I_0_11_add_573_12_lut (.I0(GND_net), .I1(n845_adj_1957[9]), 
            .I2(n576), .I3(n16520), .O(n844[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_12 (.CI(n16520), .I0(n845_adj_1957[9]), 
            .I1(n576), .CO(n16521));
    SB_LUT4 Q_15__I_0_11_add_573_11_lut (.I0(GND_net), .I1(n845_adj_1957[8]), 
            .I2(n527), .I3(n16519), .O(n844[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_11 (.CI(n16519), .I0(n845_adj_1957[8]), 
            .I1(n527), .CO(n16520));
    SB_LUT4 Q_15__I_0_i136_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n200_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i202_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n298));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i235_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n347));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_573_10_lut (.I0(GND_net), .I1(n845_adj_1957[7]), 
            .I2(n478), .I3(n16518), .O(n844[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i301_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i301_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i334_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n494));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i334_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_573_10 (.CI(n16518), .I0(n845_adj_1957[7]), 
            .I1(n478), .CO(n16519));
    SB_LUT4 Q_15__I_0_11_add_573_9_lut (.I0(GND_net), .I1(n845_adj_1957[6]), 
            .I2(n429_c), .I3(n16517), .O(n844[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_9 (.CI(n16517), .I0(n845_adj_1957[6]), 
            .I1(n429_c), .CO(n16518));
    SB_LUT4 Q_15__I_0_11_add_573_8_lut (.I0(GND_net), .I1(n845_adj_1957[5]), 
            .I2(n380), .I3(n16516), .O(n844[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_8 (.CI(n16516), .I0(n845_adj_1957[5]), 
            .I1(n380), .CO(n16517));
    SB_LUT4 Q_15__I_0_11_add_573_7_lut (.I0(GND_net), .I1(n845_adj_1957[4]), 
            .I2(n331), .I3(n16515), .O(n844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_7 (.CI(n16515), .I0(n845_adj_1957[4]), 
            .I1(n331), .CO(n16516));
    SB_LUT4 Q_15__I_0_11_add_573_6_lut (.I0(GND_net), .I1(n845_adj_1957[3]), 
            .I2(n282_c), .I3(n16514), .O(n844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_6 (.CI(n16514), .I0(n845_adj_1957[3]), 
            .I1(n282_c), .CO(n16515));
    SB_LUT4 Q_15__I_0_11_add_573_5_lut (.I0(GND_net), .I1(n845_adj_1957[2]), 
            .I2(n233_c), .I3(n16513), .O(n844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_5 (.CI(n16513), .I0(n845_adj_1957[2]), 
            .I1(n233_c), .CO(n16514));
    SB_LUT4 Q_15__I_0_11_add_573_4_lut (.I0(GND_net), .I1(n845_adj_1957[1]), 
            .I2(n184), .I3(n16512), .O(n844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_4 (.CI(n16512), .I0(n845_adj_1957[1]), 
            .I1(n184), .CO(n16513));
    SB_LUT4 Q_15__I_0_11_add_573_3_lut (.I0(GND_net), .I1(n845_adj_1957[0]), 
            .I2(n135_c), .I3(n16511), .O(n844[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_573_3 (.CI(n16511), .I0(n845_adj_1957[0]), 
            .I1(n135_c), .CO(n16512));
    SB_LUT4 Q_15__I_0_11_add_573_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n844[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_9 (.CI(n16637), .I0(n837_adj_1955[6]), 
            .I1(n429_c), .CO(n16638));
    SB_LUT4 Q_15__I_0_11_add_565_8_lut (.I0(GND_net), .I1(n837_adj_1955[5]), 
            .I2(n380), .I3(n16636), .O(n836[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_8 (.CI(n16636), .I0(n837_adj_1955[5]), 
            .I1(n380), .CO(n16637));
    SB_CARRY D_15__I_0_10_add_571_12 (.CI(n16744), .I0(n843_adj_1956[9]), 
            .I1(n570_c), .CO(n16745));
    SB_CARRY Q_15__I_0_11_add_573_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16511));
    SB_LUT4 Q_15__I_0_11_add_574_16_lut (.I0(GND_net), .I1(n846_adj_1958[13]), 
            .I2(n793), .I3(n16509), .O(n845_adj_1957[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_16 (.CI(n16509), .I0(n846_adj_1958[13]), 
            .I1(n793), .CO(n791));
    SB_LUT4 Q_15__I_0_i433_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n641));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i433_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i466_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n690));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i466_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_574_15_lut (.I0(GND_net), .I1(n846_adj_1958[12]), 
            .I2(n723), .I3(n16508), .O(n845_adj_1957[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_15 (.CI(n16508), .I0(n846_adj_1958[12]), 
            .I1(n723), .CO(n16509));
    SB_LUT4 Q_15__I_0_11_add_574_14_lut (.I0(GND_net), .I1(n846_adj_1958[11]), 
            .I2(n674), .I3(n16507), .O(n845_adj_1957[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_14 (.CI(n16507), .I0(n846_adj_1958[11]), 
            .I1(n674), .CO(n16508));
    SB_LUT4 Q_15__I_0_11_add_574_13_lut (.I0(GND_net), .I1(n846_adj_1958[10]), 
            .I2(n625_c), .I3(n16506), .O(n845_adj_1957[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_13 (.CI(n16506), .I0(n846_adj_1958[10]), 
            .I1(n625_c), .CO(n16507));
    SB_LUT4 Q_15__I_0_11_add_574_12_lut (.I0(GND_net), .I1(n846_adj_1958[9]), 
            .I2(n576), .I3(n16505), .O(n845_adj_1957[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_12 (.CI(n16505), .I0(n846_adj_1958[9]), 
            .I1(n576), .CO(n16506));
    SB_LUT4 Q_15__I_0_11_add_574_11_lut (.I0(GND_net), .I1(n846_adj_1958[8]), 
            .I2(n527), .I3(n16504), .O(n845_adj_1957[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_11 (.CI(n16504), .I0(n846_adj_1958[8]), 
            .I1(n527), .CO(n16505));
    SB_LUT4 Q_15__I_0_11_add_574_10_lut (.I0(GND_net), .I1(n846_adj_1958[7]), 
            .I2(n478), .I3(n16503), .O(n845_adj_1957[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_10 (.CI(n16503), .I0(n846_adj_1958[7]), 
            .I1(n478), .CO(n16504));
    SB_LUT4 Q_15__I_0_11_add_574_9_lut (.I0(GND_net), .I1(n846_adj_1958[6]), 
            .I2(n429_c), .I3(n16502), .O(n845_adj_1957[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_9 (.CI(n16502), .I0(n846_adj_1958[6]), 
            .I1(n429_c), .CO(n16503));
    SB_LUT4 Q_15__I_0_11_add_574_8_lut (.I0(GND_net), .I1(n846_adj_1958[5]), 
            .I2(n380), .I3(n16501), .O(n845_adj_1957[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_8 (.CI(n16501), .I0(n846_adj_1958[5]), 
            .I1(n380), .CO(n16502));
    SB_LUT4 Q_15__I_0_11_add_574_7_lut (.I0(GND_net), .I1(n846_adj_1958[4]), 
            .I2(n331), .I3(n16500), .O(n845_adj_1957[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_7 (.CI(n16500), .I0(n846_adj_1958[4]), 
            .I1(n331), .CO(n16501));
    SB_LUT4 Q_15__I_0_11_add_574_6_lut (.I0(GND_net), .I1(n846_adj_1958[3]), 
            .I2(n282_c), .I3(n16499), .O(n845_adj_1957[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_7_lut (.I0(GND_net), .I1(n837_adj_1955[4]), 
            .I2(n331), .I3(n16635), .O(n836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_6 (.CI(n16499), .I0(n846_adj_1958[3]), 
            .I1(n282_c), .CO(n16500));
    SB_LUT4 Q_15__I_0_11_add_574_5_lut (.I0(GND_net), .I1(n846_adj_1958[2]), 
            .I2(n233_c), .I3(n16498), .O(n845_adj_1957[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_5 (.CI(n16498), .I0(n846_adj_1958[2]), 
            .I1(n233_c), .CO(n16499));
    SB_LUT4 Q_15__I_0_11_add_574_4_lut (.I0(GND_net), .I1(n846_adj_1958[1]), 
            .I2(n184), .I3(n16497), .O(n845_adj_1957[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_7 (.CI(n16635), .I0(n837_adj_1955[4]), 
            .I1(n331), .CO(n16636));
    SB_CARRY Q_15__I_0_11_add_574_4 (.CI(n16497), .I0(n846_adj_1958[1]), 
            .I1(n184), .CO(n16498));
    SB_LUT4 Q_15__I_0_11_add_574_3_lut (.I0(GND_net), .I1(n846_adj_1958[0]), 
            .I2(n135_c), .I3(n16496), .O(n845_adj_1957[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_3 (.CI(n16496), .I0(n846_adj_1958[0]), 
            .I1(n135_c), .CO(n16497));
    SB_LUT4 Q_15__I_0_11_add_574_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n845_adj_1957[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_574_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16496));
    SB_LUT4 Q_15__I_0_11_add_575_16_lut (.I0(GND_net), .I1(n19680), .I2(n793), 
            .I3(n16495), .O(n846_adj_1958[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_575_15_lut (.I0(GND_net), .I1(n685_adj_1082), 
            .I2(n723), .I3(n16494), .O(n846_adj_1958[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_15 (.CI(n16494), .I0(n685_adj_1082), .I1(n723), 
            .CO(n16495));
    SB_LUT4 Q_15__I_0_11_add_575_14_lut (.I0(GND_net), .I1(n636_adj_1083), 
            .I2(n674), .I3(n16493), .O(n846_adj_1958[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_14 (.CI(n16493), .I0(n636_adj_1083), .I1(n674), 
            .CO(n16494));
    SB_LUT4 Q_15__I_0_11_add_575_13_lut (.I0(GND_net), .I1(n587_adj_203), 
            .I2(n625_c), .I3(n16492), .O(n846_adj_1958[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_13 (.CI(n16492), .I0(n587_adj_203), .I1(n625_c), 
            .CO(n16493));
    SB_LUT4 Q_15__I_0_11_add_575_12_lut (.I0(GND_net), .I1(n538_c), .I2(n576), 
            .I3(n16491), .O(n846_adj_1958[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_12 (.CI(n16491), .I0(n538_c), .I1(n576), 
            .CO(n16492));
    SB_LUT4 Q_15__I_0_11_add_575_11_lut (.I0(GND_net), .I1(n489), .I2(n527), 
            .I3(n16490), .O(n846_adj_1958[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_11 (.CI(n16490), .I0(n489), .I1(n527), 
            .CO(n16491));
    SB_LUT4 Q_15__I_0_11_add_575_10_lut (.I0(GND_net), .I1(n440), .I2(n478), 
            .I3(n16489), .O(n846_adj_1958[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_10 (.CI(n16489), .I0(n440), .I1(n478), 
            .CO(n16490));
    SB_LUT4 Q_15__I_0_11_add_575_9_lut (.I0(GND_net), .I1(n391), .I2(n429_c), 
            .I3(n16488), .O(n846_adj_1958[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_9 (.CI(n16488), .I0(n391), .I1(n429_c), 
            .CO(n16489));
    SB_LUT4 Q_15__I_0_11_add_575_8_lut (.I0(GND_net), .I1(n342), .I2(n380), 
            .I3(n16487), .O(n846_adj_1958[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_8 (.CI(n16487), .I0(n342), .I1(n380), 
            .CO(n16488));
    SB_LUT4 Q_15__I_0_11_add_565_6_lut (.I0(GND_net), .I1(n837_adj_1955[3]), 
            .I2(n282_c), .I3(n16634), .O(n836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_6 (.CI(n16634), .I0(n837_adj_1955[3]), 
            .I1(n282_c), .CO(n16635));
    SB_LUT4 Q_15__I_0_11_add_575_7_lut (.I0(GND_net), .I1(n293), .I2(n331), 
            .I3(n16486), .O(n846_adj_1958[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_7 (.CI(n16486), .I0(n293), .I1(n331), 
            .CO(n16487));
    SB_LUT4 Q_15__I_0_11_add_565_5_lut (.I0(GND_net), .I1(n837_adj_1955[2]), 
            .I2(n233_c), .I3(n16633), .O(n836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_575_6_lut (.I0(GND_net), .I1(n244_c), .I2(n282_c), 
            .I3(n16485), .O(n846_adj_1958[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_6 (.CI(n16485), .I0(n244_c), .I1(n282_c), 
            .CO(n16486));
    SB_LUT4 Q_15__I_0_11_add_575_5_lut (.I0(GND_net), .I1(n195_c), .I2(n233_c), 
            .I3(n16484), .O(n846_adj_1958[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_5 (.CI(n16484), .I0(n195_c), .I1(n233_c), 
            .CO(n16485));
    SB_LUT4 Q_15__I_0_11_add_575_4_lut (.I0(GND_net), .I1(n146), .I2(n184), 
            .I3(n16483), .O(n846_adj_1958[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_4 (.CI(n16483), .I0(n146), .I1(n184), 
            .CO(n16484));
    SB_LUT4 Q_15__I_0_11_add_575_3_lut (.I0(GND_net), .I1(n97), .I2(n135_c), 
            .I3(n16482), .O(n846_adj_1958[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_3 (.CI(n16482), .I0(n97), .I1(n135_c), 
            .CO(n16483));
    SB_LUT4 Q_15__I_0_11_add_575_2_lut (.I0(GND_net), .I1(n48), .I2(n86), 
            .I3(GND_net), .O(n846_adj_1958[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_575_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_575_2 (.CI(GND_net), .I0(n48), .I1(n86), 
            .CO(n16482));
    SB_LUT4 add_1230_16_lut (.I0(GND_net), .I1(n846[14]), .I2(n791_adj_1086), 
            .I3(n16481), .O(Product1_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1230_15_lut (.I0(GND_net), .I1(n845[14]), .I2(n787_adj_1088), 
            .I3(n16480), .O(Product1_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_15 (.CI(n16480), .I0(n845[14]), .I1(n787_adj_1088), 
            .CO(n16481));
    SB_LUT4 add_1230_14_lut (.I0(GND_net), .I1(n844_adj_1959[14]), .I2(n783_adj_1090), 
            .I3(n16479), .O(Product1_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_14 (.CI(n16479), .I0(n844_adj_1959[14]), .I1(n783_adj_1090), 
            .CO(n16480));
    SB_LUT4 add_1230_13_lut (.I0(GND_net), .I1(n843_adj_1956[14]), .I2(n779_adj_1067), 
            .I3(n16478), .O(Product1_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_13 (.CI(n16478), .I0(n843_adj_1956[14]), .I1(n779_adj_1067), 
            .CO(n16479));
    SB_LUT4 add_1230_12_lut (.I0(GND_net), .I1(n842_adj_1954[14]), .I2(n775), 
            .I3(n16477), .O(Product1_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_12 (.CI(n16477), .I0(n842_adj_1954[14]), .I1(n775), 
            .CO(n16478));
    SB_LUT4 add_1230_11_lut (.I0(GND_net), .I1(n841[14]), .I2(n771), .I3(n16476), 
            .O(Product1_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_11 (.CI(n16476), .I0(n841[14]), .I1(n771), .CO(n16477));
    SB_LUT4 add_1230_10_lut (.I0(GND_net), .I1(n840_adj_1950[14]), .I2(n767_adj_1092), 
            .I3(n16475), .O(Product1_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_10 (.CI(n16475), .I0(n840_adj_1950[14]), .I1(n767_adj_1092), 
            .CO(n16476));
    SB_LUT4 add_1230_9_lut (.I0(GND_net), .I1(n839_adj_1951[14]), .I2(n763), 
            .I3(n16474), .O(Product1_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_9 (.CI(n16474), .I0(n839_adj_1951[14]), .I1(n763), 
            .CO(n16475));
    SB_LUT4 add_1230_8_lut (.I0(GND_net), .I1(n838[14]), .I2(n759), .I3(n16473), 
            .O(Product1_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_8 (.CI(n16473), .I0(n838[14]), .I1(n759), .CO(n16474));
    SB_LUT4 add_1230_7_lut (.I0(GND_net), .I1(n837[14]), .I2(n755_adj_1094), 
            .I3(n16472), .O(Product1_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_7 (.CI(n16472), .I0(n837[14]), .I1(n755_adj_1094), 
            .CO(n16473));
    SB_LUT4 add_1230_6_lut (.I0(GND_net), .I1(n836_adj_1960[14]), .I2(n751), 
            .I3(n16471), .O(Product1_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_6 (.CI(n16471), .I0(n836_adj_1960[14]), .I1(n751), 
            .CO(n16472));
    SB_LUT4 add_1230_5_lut (.I0(GND_net), .I1(n835_adj_1961[14]), .I2(n747), 
            .I3(n16470), .O(Product1_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_11_lut (.I0(GND_net), .I1(n843_adj_1956[8]), 
            .I2(n521), .I3(n16743), .O(n842_adj_1954[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_5 (.CI(n16470), .I0(n835_adj_1961[14]), .I1(n747), 
            .CO(n16471));
    SB_LUT4 add_1230_4_lut (.I0(GND_net), .I1(n834[14]), .I2(n743), .I3(n16469), 
            .O(Product1_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_4 (.CI(n16469), .I0(n834[14]), .I1(n743), .CO(n16470));
    SB_LUT4 add_1230_3_lut (.I0(GND_net), .I1(n833[14]), .I2(n739), .I3(n16468), 
            .O(Product1_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_5 (.CI(n16633), .I0(n837_adj_1955[2]), 
            .I1(n233_c), .CO(n16634));
    SB_CARRY D_15__I_0_10_add_571_11 (.CI(n16743), .I0(n843_adj_1956[8]), 
            .I1(n521), .CO(n16744));
    SB_CARRY add_1230_3 (.CI(n16468), .I0(n833[14]), .I1(n739), .CO(n16469));
    SB_LUT4 add_1230_2_lut (.I0(GND_net), .I1(\dVoltage[15] ), .I2(Look_Up_Table_out1_1[15]), 
            .I3(n16467), .O(Product1_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1230_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1230_2 (.CI(n16467), .I0(\dVoltage[15] ), .I1(Look_Up_Table_out1_1[15]), 
            .CO(n16468));
    SB_CARRY add_1230_1 (.CI(GND_net), .I0(n832[14]), .I1(n832[14]), .CO(n16467));
    SB_LUT4 D_15__I_0_add_563_16_lut (.I0(GND_net), .I1(n835_adj_1963[13]), 
            .I2(n793_adj_1098), .I3(n16465), .O(n834_adj_1962[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_16 (.CI(n16465), .I0(n835_adj_1963[13]), 
            .I1(n793_adj_1098), .CO(n747_adj_1099));
    SB_LUT4 D_15__I_0_add_563_15_lut (.I0(GND_net), .I1(n835_adj_1963[12]), 
            .I2(n723_adj_1100), .I3(n16464), .O(n834_adj_1962[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_15 (.CI(n16464), .I0(n835_adj_1963[12]), 
            .I1(n723_adj_1100), .CO(n16465));
    SB_LUT4 D_15__I_0_add_563_14_lut (.I0(GND_net), .I1(n835_adj_1963[11]), 
            .I2(n674_adj_1101), .I3(n16463), .O(n833_adj_1964[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_14 (.CI(n16463), .I0(n835_adj_1963[11]), 
            .I1(n674_adj_1101), .CO(n16464));
    SB_LUT4 D_15__I_0_add_563_13_lut (.I0(GND_net), .I1(n835_adj_1963[10]), 
            .I2(n625_adj_1102), .I3(n16462), .O(Product3_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_13 (.CI(n16462), .I0(n835_adj_1963[10]), 
            .I1(n625_adj_1102), .CO(n16463));
    SB_LUT4 D_15__I_0_add_563_12_lut (.I0(GND_net), .I1(n835_adj_1963[9]), 
            .I2(n576_adj_1104), .I3(n16461), .O(Product3_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_12 (.CI(n16461), .I0(n835_adj_1963[9]), .I1(n576_adj_1104), 
            .CO(n16462));
    SB_LUT4 D_15__I_0_add_563_11_lut (.I0(GND_net), .I1(n835_adj_1963[8]), 
            .I2(n527_adj_1106), .I3(n16460), .O(Product3_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_11 (.CI(n16460), .I0(n835_adj_1963[8]), .I1(n527_adj_1106), 
            .CO(n16461));
    SB_LUT4 D_15__I_0_add_563_10_lut (.I0(GND_net), .I1(n835_adj_1963[7]), 
            .I2(n478_adj_1108), .I3(n16459), .O(Product3_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_10 (.CI(n16459), .I0(n835_adj_1963[7]), .I1(n478_adj_1108), 
            .CO(n16460));
    SB_LUT4 D_15__I_0_add_563_9_lut (.I0(GND_net), .I1(n835_adj_1963[6]), 
            .I2(n429_adj_1110), .I3(n16458), .O(Product3_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_9 (.CI(n16458), .I0(n835_adj_1963[6]), .I1(n429_adj_1110), 
            .CO(n16459));
    SB_LUT4 D_15__I_0_add_563_8_lut (.I0(GND_net), .I1(n835_adj_1963[5]), 
            .I2(n380_adj_1112), .I3(n16457), .O(Product3_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_8 (.CI(n16457), .I0(n835_adj_1963[5]), .I1(n380_adj_1112), 
            .CO(n16458));
    SB_LUT4 D_15__I_0_add_563_7_lut (.I0(GND_net), .I1(n835_adj_1963[4]), 
            .I2(n331_adj_1114), .I3(n16456), .O(Product3_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_7 (.CI(n16456), .I0(n835_adj_1963[4]), .I1(n331_adj_1114), 
            .CO(n16457));
    SB_LUT4 D_15__I_0_add_563_6_lut (.I0(GND_net), .I1(n835_adj_1963[3]), 
            .I2(n282_adj_1116), .I3(n16455), .O(Product3_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_6 (.CI(n16455), .I0(n835_adj_1963[3]), .I1(n282_adj_1116), 
            .CO(n16456));
    SB_LUT4 D_15__I_0_add_563_5_lut (.I0(GND_net), .I1(n835_adj_1963[2]), 
            .I2(n233), .I3(n16454), .O(Product3_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_5 (.CI(n16454), .I0(n835_adj_1963[2]), .I1(n233), 
            .CO(n16455));
    SB_LUT4 D_15__I_0_add_563_4_lut (.I0(GND_net), .I1(n835_adj_1963[1]), 
            .I2(n184_adj_1120), .I3(n16453), .O(Product3_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_4_lut (.I0(GND_net), .I1(n837_adj_1955[1]), 
            .I2(n184), .I3(n16632), .O(n836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_4 (.CI(n16453), .I0(n835_adj_1963[1]), .I1(n184_adj_1120), 
            .CO(n16454));
    SB_LUT4 D_15__I_0_add_563_3_lut (.I0(GND_net), .I1(n835_adj_1963[0]), 
            .I2(n135_adj_1123), .I3(n16452), .O(Product3_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_3 (.CI(n16452), .I0(n835_adj_1963[0]), .I1(n135_adj_1123), 
            .CO(n16453));
    SB_LUT4 D_15__I_0_add_563_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(Product3_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_563_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16452));
    SB_LUT4 D_15__I_0_add_564_16_lut (.I0(GND_net), .I1(n836_adj_1965[13]), 
            .I2(n793_adj_1098), .I3(n16450), .O(n835_adj_1963[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_16 (.CI(n16450), .I0(n836_adj_1965[13]), 
            .I1(n793_adj_1098), .CO(n751_adj_1127));
    SB_LUT4 D_15__I_0_add_564_15_lut (.I0(GND_net), .I1(n836_adj_1965[12]), 
            .I2(n723_adj_1100), .I3(n16449), .O(n835_adj_1963[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_15 (.CI(n16449), .I0(n836_adj_1965[12]), 
            .I1(n723_adj_1100), .CO(n16450));
    SB_LUT4 D_15__I_0_add_564_14_lut (.I0(GND_net), .I1(n836_adj_1965[11]), 
            .I2(n674_adj_1101), .I3(n16448), .O(n835_adj_1963[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_14 (.CI(n16448), .I0(n836_adj_1965[11]), 
            .I1(n674_adj_1101), .CO(n16449));
    SB_LUT4 D_15__I_0_add_564_13_lut (.I0(GND_net), .I1(n836_adj_1965[10]), 
            .I2(n625_adj_1102), .I3(n16447), .O(n835_adj_1963[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_565_4 (.CI(n16632), .I0(n837_adj_1955[1]), 
            .I1(n184), .CO(n16633));
    SB_LUT4 D_15__I_0_10_add_571_10_lut (.I0(GND_net), .I1(n843_adj_1956[7]), 
            .I2(n472), .I3(n16742), .O(n842_adj_1954[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_13 (.CI(n16447), .I0(n836_adj_1965[10]), 
            .I1(n625_adj_1102), .CO(n16448));
    SB_LUT4 D_15__I_0_add_564_12_lut (.I0(GND_net), .I1(n836_adj_1965[9]), 
            .I2(n576_adj_1104), .I3(n16446), .O(n835_adj_1963[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_12 (.CI(n16446), .I0(n836_adj_1965[9]), .I1(n576_adj_1104), 
            .CO(n16447));
    SB_LUT4 D_15__I_0_add_564_11_lut (.I0(GND_net), .I1(n836_adj_1965[8]), 
            .I2(n527_adj_1106), .I3(n16445), .O(n835_adj_1963[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_11 (.CI(n16445), .I0(n836_adj_1965[8]), .I1(n527_adj_1106), 
            .CO(n16446));
    SB_LUT4 D_15__I_0_add_564_10_lut (.I0(GND_net), .I1(n836_adj_1965[7]), 
            .I2(n478_adj_1108), .I3(n16444), .O(n835_adj_1963[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_10 (.CI(n16444), .I0(n836_adj_1965[7]), .I1(n478_adj_1108), 
            .CO(n16445));
    SB_LUT4 D_15__I_0_add_564_9_lut (.I0(GND_net), .I1(n836_adj_1965[6]), 
            .I2(n429_adj_1110), .I3(n16443), .O(n835_adj_1963[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_9 (.CI(n16443), .I0(n836_adj_1965[6]), .I1(n429_adj_1110), 
            .CO(n16444));
    SB_LUT4 D_15__I_0_add_564_8_lut (.I0(GND_net), .I1(n836_adj_1965[5]), 
            .I2(n380_adj_1112), .I3(n16442), .O(n835_adj_1963[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_8 (.CI(n16442), .I0(n836_adj_1965[5]), .I1(n380_adj_1112), 
            .CO(n16443));
    SB_LUT4 D_15__I_0_add_564_7_lut (.I0(GND_net), .I1(n836_adj_1965[4]), 
            .I2(n331_adj_1114), .I3(n16441), .O(n835_adj_1963[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_7 (.CI(n16441), .I0(n836_adj_1965[4]), .I1(n331_adj_1114), 
            .CO(n16442));
    SB_LUT4 D_15__I_0_add_564_6_lut (.I0(GND_net), .I1(n836_adj_1965[3]), 
            .I2(n282_adj_1116), .I3(n16440), .O(n835_adj_1963[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_6 (.CI(n16440), .I0(n836_adj_1965[3]), .I1(n282_adj_1116), 
            .CO(n16441));
    SB_LUT4 D_15__I_0_add_564_5_lut (.I0(GND_net), .I1(n836_adj_1965[2]), 
            .I2(n233), .I3(n16439), .O(n835_adj_1963[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_5 (.CI(n16439), .I0(n836_adj_1965[2]), .I1(n233), 
            .CO(n16440));
    SB_LUT4 D_15__I_0_add_564_4_lut (.I0(GND_net), .I1(n836_adj_1965[1]), 
            .I2(n184_adj_1120), .I3(n16438), .O(n835_adj_1963[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_4 (.CI(n16438), .I0(n836_adj_1965[1]), .I1(n184_adj_1120), 
            .CO(n16439));
    SB_LUT4 D_15__I_0_add_564_3_lut (.I0(GND_net), .I1(n836_adj_1965[0]), 
            .I2(n135_adj_1123), .I3(n16437), .O(n835_adj_1963[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_3 (.CI(n16437), .I0(n836_adj_1965[0]), .I1(n135_adj_1123), 
            .CO(n16438));
    SB_LUT4 D_15__I_0_add_564_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n835_adj_1963[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_564_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16437));
    SB_LUT4 D_15__I_0_add_565_16_lut (.I0(GND_net), .I1(n837_adj_1966[13]), 
            .I2(n793_adj_1098), .I3(n16435), .O(n836_adj_1965[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_16 (.CI(n16435), .I0(n837_adj_1966[13]), 
            .I1(n793_adj_1098), .CO(n755_adj_1144));
    SB_LUT4 D_15__I_0_add_565_15_lut (.I0(GND_net), .I1(n837_adj_1966[12]), 
            .I2(n723_adj_1100), .I3(n16434), .O(n836_adj_1965[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_15 (.CI(n16434), .I0(n837_adj_1966[12]), 
            .I1(n723_adj_1100), .CO(n16435));
    SB_LUT4 D_15__I_0_add_565_14_lut (.I0(GND_net), .I1(n837_adj_1966[11]), 
            .I2(n674_adj_1101), .I3(n16433), .O(n836_adj_1965[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_14 (.CI(n16433), .I0(n837_adj_1966[11]), 
            .I1(n674_adj_1101), .CO(n16434));
    SB_LUT4 D_15__I_0_add_565_13_lut (.I0(GND_net), .I1(n837_adj_1966[10]), 
            .I2(n625_adj_1102), .I3(n16432), .O(n836_adj_1965[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_13 (.CI(n16432), .I0(n837_adj_1966[10]), 
            .I1(n625_adj_1102), .CO(n16433));
    SB_LUT4 D_15__I_0_add_565_12_lut (.I0(GND_net), .I1(n837_adj_1966[9]), 
            .I2(n576_adj_1104), .I3(n16431), .O(n836_adj_1965[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_12 (.CI(n16431), .I0(n837_adj_1966[9]), .I1(n576_adj_1104), 
            .CO(n16432));
    SB_LUT4 D_15__I_0_add_565_11_lut (.I0(GND_net), .I1(n837_adj_1966[8]), 
            .I2(n527_adj_1106), .I3(n16430), .O(n836_adj_1965[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_11 (.CI(n16430), .I0(n837_adj_1966[8]), .I1(n527_adj_1106), 
            .CO(n16431));
    SB_LUT4 D_15__I_0_add_565_10_lut (.I0(GND_net), .I1(n837_adj_1966[7]), 
            .I2(n478_adj_1108), .I3(n16429), .O(n836_adj_1965[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_10 (.CI(n16429), .I0(n837_adj_1966[7]), .I1(n478_adj_1108), 
            .CO(n16430));
    SB_LUT4 D_15__I_0_add_565_9_lut (.I0(GND_net), .I1(n837_adj_1966[6]), 
            .I2(n429_adj_1110), .I3(n16428), .O(n836_adj_1965[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_9 (.CI(n16428), .I0(n837_adj_1966[6]), .I1(n429_adj_1110), 
            .CO(n16429));
    SB_LUT4 D_15__I_0_add_565_8_lut (.I0(GND_net), .I1(n837_adj_1966[5]), 
            .I2(n380_adj_1112), .I3(n16427), .O(n836_adj_1965[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_8 (.CI(n16427), .I0(n837_adj_1966[5]), .I1(n380_adj_1112), 
            .CO(n16428));
    SB_LUT4 D_15__I_0_add_565_7_lut (.I0(GND_net), .I1(n837_adj_1966[4]), 
            .I2(n331_adj_1114), .I3(n16426), .O(n836_adj_1965[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_7 (.CI(n16426), .I0(n837_adj_1966[4]), .I1(n331_adj_1114), 
            .CO(n16427));
    SB_LUT4 D_15__I_0_add_565_6_lut (.I0(GND_net), .I1(n837_adj_1966[3]), 
            .I2(n282_adj_1116), .I3(n16425), .O(n836_adj_1965[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_6 (.CI(n16425), .I0(n837_adj_1966[3]), .I1(n282_adj_1116), 
            .CO(n16426));
    SB_LUT4 D_15__I_0_add_565_5_lut (.I0(GND_net), .I1(n837_adj_1966[2]), 
            .I2(n233), .I3(n16424), .O(n836_adj_1965[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_5 (.CI(n16424), .I0(n837_adj_1966[2]), .I1(n233), 
            .CO(n16425));
    SB_LUT4 D_15__I_0_add_565_4_lut (.I0(GND_net), .I1(n837_adj_1966[1]), 
            .I2(n184_adj_1120), .I3(n16423), .O(n836_adj_1965[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_4 (.CI(n16423), .I0(n837_adj_1966[1]), .I1(n184_adj_1120), 
            .CO(n16424));
    SB_LUT4 D_15__I_0_add_565_3_lut (.I0(GND_net), .I1(n837_adj_1966[0]), 
            .I2(n135_adj_1123), .I3(n16422), .O(n836_adj_1965[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_3 (.CI(n16422), .I0(n837_adj_1966[0]), .I1(n135_adj_1123), 
            .CO(n16423));
    SB_LUT4 D_15__I_0_add_565_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n836_adj_1965[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_565_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16422));
    SB_LUT4 D_15__I_0_add_566_16_lut (.I0(GND_net), .I1(n838_adj_1967[13]), 
            .I2(n793_adj_1098), .I3(n16420), .O(n837_adj_1966[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_16 (.CI(n16420), .I0(n838_adj_1967[13]), 
            .I1(n793_adj_1098), .CO(n759_adj_1158));
    SB_LUT4 D_15__I_0_add_566_15_lut (.I0(GND_net), .I1(n838_adj_1967[12]), 
            .I2(n723_adj_1100), .I3(n16419), .O(n837_adj_1966[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_15 (.CI(n16419), .I0(n838_adj_1967[12]), 
            .I1(n723_adj_1100), .CO(n16420));
    SB_LUT4 D_15__I_0_add_566_14_lut (.I0(GND_net), .I1(n838_adj_1967[11]), 
            .I2(n674_adj_1101), .I3(n16418), .O(n837_adj_1966[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_14 (.CI(n16418), .I0(n838_adj_1967[11]), 
            .I1(n674_adj_1101), .CO(n16419));
    SB_LUT4 D_15__I_0_add_566_13_lut (.I0(GND_net), .I1(n838_adj_1967[10]), 
            .I2(n625_adj_1102), .I3(n16417), .O(n837_adj_1966[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_13 (.CI(n16417), .I0(n838_adj_1967[10]), 
            .I1(n625_adj_1102), .CO(n16418));
    SB_LUT4 D_15__I_0_add_566_12_lut (.I0(GND_net), .I1(n838_adj_1967[9]), 
            .I2(n576_adj_1104), .I3(n16416), .O(n837_adj_1966[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_12 (.CI(n16416), .I0(n838_adj_1967[9]), .I1(n576_adj_1104), 
            .CO(n16417));
    SB_LUT4 D_15__I_0_add_566_11_lut (.I0(GND_net), .I1(n838_adj_1967[8]), 
            .I2(n527_adj_1106), .I3(n16415), .O(n837_adj_1966[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_11 (.CI(n16415), .I0(n838_adj_1967[8]), .I1(n527_adj_1106), 
            .CO(n16416));
    SB_LUT4 D_15__I_0_add_566_10_lut (.I0(GND_net), .I1(n838_adj_1967[7]), 
            .I2(n478_adj_1108), .I3(n16414), .O(n837_adj_1966[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_10 (.CI(n16414), .I0(n838_adj_1967[7]), .I1(n478_adj_1108), 
            .CO(n16415));
    SB_LUT4 D_15__I_0_add_566_9_lut (.I0(GND_net), .I1(n838_adj_1967[6]), 
            .I2(n429_adj_1110), .I3(n16413), .O(n837_adj_1966[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_9 (.CI(n16413), .I0(n838_adj_1967[6]), .I1(n429_adj_1110), 
            .CO(n16414));
    SB_LUT4 D_15__I_0_add_566_8_lut (.I0(GND_net), .I1(n838_adj_1967[5]), 
            .I2(n380_adj_1112), .I3(n16412), .O(n837_adj_1966[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_8 (.CI(n16412), .I0(n838_adj_1967[5]), .I1(n380_adj_1112), 
            .CO(n16413));
    SB_LUT4 D_15__I_0_add_566_7_lut (.I0(GND_net), .I1(n838_adj_1967[4]), 
            .I2(n331_adj_1114), .I3(n16411), .O(n837_adj_1966[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_7 (.CI(n16411), .I0(n838_adj_1967[4]), .I1(n331_adj_1114), 
            .CO(n16412));
    SB_LUT4 D_15__I_0_add_566_6_lut (.I0(GND_net), .I1(n838_adj_1967[3]), 
            .I2(n282_adj_1116), .I3(n16410), .O(n837_adj_1966[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_6 (.CI(n16410), .I0(n838_adj_1967[3]), .I1(n282_adj_1116), 
            .CO(n16411));
    SB_LUT4 D_15__I_0_add_566_5_lut (.I0(GND_net), .I1(n838_adj_1967[2]), 
            .I2(n233), .I3(n16409), .O(n837_adj_1966[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_3_lut (.I0(GND_net), .I1(n837_adj_1955[0]), 
            .I2(n135_c), .I3(n16631), .O(n836[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_5 (.CI(n16409), .I0(n838_adj_1967[2]), .I1(n233), 
            .CO(n16410));
    SB_LUT4 D_15__I_0_add_566_4_lut (.I0(GND_net), .I1(n838_adj_1967[1]), 
            .I2(n184_adj_1120), .I3(n16408), .O(n837_adj_1966[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_10 (.CI(n16742), .I0(n843_adj_1956[7]), 
            .I1(n472), .CO(n16743));
    SB_CARRY D_15__I_0_add_566_4 (.CI(n16408), .I0(n838_adj_1967[1]), .I1(n184_adj_1120), 
            .CO(n16409));
    SB_LUT4 D_15__I_0_add_566_3_lut (.I0(GND_net), .I1(n838_adj_1967[0]), 
            .I2(n135_adj_1123), .I3(n16407), .O(n837_adj_1966[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_3 (.CI(n16407), .I0(n838_adj_1967[0]), .I1(n135_adj_1123), 
            .CO(n16408));
    SB_LUT4 D_15__I_0_add_566_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n837_adj_1966[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_566_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16407));
    SB_LUT4 D_15__I_0_add_567_16_lut (.I0(GND_net), .I1(n839_adj_1968[13]), 
            .I2(n793_adj_1098), .I3(n16405), .O(n838_adj_1967[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_16 (.CI(n16405), .I0(n839_adj_1968[13]), 
            .I1(n793_adj_1098), .CO(n763_adj_1175));
    SB_LUT4 D_15__I_0_add_567_15_lut (.I0(GND_net), .I1(n839_adj_1968[12]), 
            .I2(n723_adj_1100), .I3(n16404), .O(n838_adj_1967[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_15 (.CI(n16404), .I0(n839_adj_1968[12]), 
            .I1(n723_adj_1100), .CO(n16405));
    SB_LUT4 D_15__I_0_add_567_14_lut (.I0(GND_net), .I1(n839_adj_1968[11]), 
            .I2(n674_adj_1101), .I3(n16403), .O(n838_adj_1967[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_14 (.CI(n16403), .I0(n839_adj_1968[11]), 
            .I1(n674_adj_1101), .CO(n16404));
    SB_LUT4 D_15__I_0_add_567_13_lut (.I0(GND_net), .I1(n839_adj_1968[10]), 
            .I2(n625_adj_1102), .I3(n16402), .O(n838_adj_1967[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_13 (.CI(n16402), .I0(n839_adj_1968[10]), 
            .I1(n625_adj_1102), .CO(n16403));
    SB_LUT4 D_15__I_0_add_567_12_lut (.I0(GND_net), .I1(n839_adj_1968[9]), 
            .I2(n576_adj_1104), .I3(n16401), .O(n838_adj_1967[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_12 (.CI(n16401), .I0(n839_adj_1968[9]), .I1(n576_adj_1104), 
            .CO(n16402));
    SB_LUT4 D_15__I_0_add_567_11_lut (.I0(GND_net), .I1(n839_adj_1968[8]), 
            .I2(n527_adj_1106), .I3(n16400), .O(n838_adj_1967[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_11 (.CI(n16400), .I0(n839_adj_1968[8]), .I1(n527_adj_1106), 
            .CO(n16401));
    SB_LUT4 D_15__I_0_add_567_10_lut (.I0(GND_net), .I1(n839_adj_1968[7]), 
            .I2(n478_adj_1108), .I3(n16399), .O(n838_adj_1967[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_10 (.CI(n16399), .I0(n839_adj_1968[7]), .I1(n478_adj_1108), 
            .CO(n16400));
    SB_LUT4 D_15__I_0_add_567_9_lut (.I0(GND_net), .I1(n839_adj_1968[6]), 
            .I2(n429_adj_1110), .I3(n16398), .O(n838_adj_1967[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_9 (.CI(n16398), .I0(n839_adj_1968[6]), .I1(n429_adj_1110), 
            .CO(n16399));
    SB_LUT4 D_15__I_0_add_567_8_lut (.I0(GND_net), .I1(n839_adj_1968[5]), 
            .I2(n380_adj_1112), .I3(n16397), .O(n838_adj_1967[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_8 (.CI(n16397), .I0(n839_adj_1968[5]), .I1(n380_adj_1112), 
            .CO(n16398));
    SB_LUT4 D_15__I_0_add_567_7_lut (.I0(GND_net), .I1(n839_adj_1968[4]), 
            .I2(n331_adj_1114), .I3(n16396), .O(n838_adj_1967[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_15 (.CI(n16598), .I0(n840[12]), .I1(n723), 
            .CO(n16599));
    SB_CARRY D_15__I_0_10_add_575_13 (.CI(n16686), .I0(n587), .I1(n631), 
            .CO(n16687));
    SB_CARRY D_15__I_0_add_567_7 (.CI(n16396), .I0(n839_adj_1968[4]), .I1(n331_adj_1114), 
            .CO(n16397));
    SB_LUT4 D_15__I_0_add_567_6_lut (.I0(GND_net), .I1(n839_adj_1968[3]), 
            .I2(n282_adj_1116), .I3(n16395), .O(n838_adj_1967[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_6 (.CI(n16395), .I0(n839_adj_1968[3]), .I1(n282_adj_1116), 
            .CO(n16396));
    SB_LUT4 D_15__I_0_add_567_5_lut (.I0(GND_net), .I1(n839_adj_1968[2]), 
            .I2(n233), .I3(n16394), .O(n838_adj_1967[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_5 (.CI(n16394), .I0(n839_adj_1968[2]), .I1(n233), 
            .CO(n16395));
    SB_LUT4 D_15__I_0_add_567_4_lut (.I0(GND_net), .I1(n839_adj_1968[1]), 
            .I2(n184_adj_1120), .I3(n16393), .O(n838_adj_1967[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_4 (.CI(n16393), .I0(n839_adj_1968[1]), .I1(n184_adj_1120), 
            .CO(n16394));
    SB_LUT4 D_15__I_0_add_567_3_lut (.I0(GND_net), .I1(n839_adj_1968[0]), 
            .I2(n135_adj_1123), .I3(n16392), .O(n838_adj_1967[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_3 (.CI(n16392), .I0(n839_adj_1968[0]), .I1(n135_adj_1123), 
            .CO(n16393));
    SB_LUT4 D_15__I_0_add_567_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n838_adj_1967[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_567_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16392));
    SB_LUT4 D_15__I_0_add_568_16_lut (.I0(GND_net), .I1(n840_adj_1969[13]), 
            .I2(n793_adj_1098), .I3(n16390), .O(n839_adj_1968[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_16 (.CI(n16390), .I0(n840_adj_1969[13]), 
            .I1(n793_adj_1098), .CO(n767_adj_1191));
    SB_LUT4 D_15__I_0_add_568_15_lut (.I0(GND_net), .I1(n840_adj_1969[12]), 
            .I2(n723_adj_1100), .I3(n16389), .O(n839_adj_1968[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_15 (.CI(n16389), .I0(n840_adj_1969[12]), 
            .I1(n723_adj_1100), .CO(n16390));
    SB_LUT4 D_15__I_0_add_568_14_lut (.I0(GND_net), .I1(n840_adj_1969[11]), 
            .I2(n674_adj_1101), .I3(n16388), .O(n839_adj_1968[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_14 (.CI(n16388), .I0(n840_adj_1969[11]), 
            .I1(n674_adj_1101), .CO(n16389));
    SB_LUT4 D_15__I_0_add_568_13_lut (.I0(GND_net), .I1(n840_adj_1969[10]), 
            .I2(n625_adj_1102), .I3(n16387), .O(n839_adj_1968[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_13 (.CI(n16387), .I0(n840_adj_1969[10]), 
            .I1(n625_adj_1102), .CO(n16388));
    SB_LUT4 D_15__I_0_add_568_12_lut (.I0(GND_net), .I1(n840_adj_1969[9]), 
            .I2(n576_adj_1104), .I3(n16386), .O(n839_adj_1968[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_12 (.CI(n16386), .I0(n840_adj_1969[9]), .I1(n576_adj_1104), 
            .CO(n16387));
    SB_LUT4 D_15__I_0_add_568_11_lut (.I0(GND_net), .I1(n840_adj_1969[8]), 
            .I2(n527_adj_1106), .I3(n16385), .O(n839_adj_1968[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_11 (.CI(n16385), .I0(n840_adj_1969[8]), .I1(n527_adj_1106), 
            .CO(n16386));
    SB_LUT4 D_15__I_0_add_568_10_lut (.I0(GND_net), .I1(n840_adj_1969[7]), 
            .I2(n478_adj_1108), .I3(n16384), .O(n839_adj_1968[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_10 (.CI(n16384), .I0(n840_adj_1969[7]), .I1(n478_adj_1108), 
            .CO(n16385));
    SB_LUT4 D_15__I_0_add_568_9_lut (.I0(GND_net), .I1(n840_adj_1969[6]), 
            .I2(n429_adj_1110), .I3(n16383), .O(n839_adj_1968[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_9 (.CI(n16383), .I0(n840_adj_1969[6]), .I1(n429_adj_1110), 
            .CO(n16384));
    SB_LUT4 D_15__I_0_add_568_8_lut (.I0(GND_net), .I1(n840_adj_1969[5]), 
            .I2(n380_adj_1112), .I3(n16382), .O(n839_adj_1968[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_8 (.CI(n16382), .I0(n840_adj_1969[5]), .I1(n380_adj_1112), 
            .CO(n16383));
    SB_LUT4 D_15__I_0_add_568_7_lut (.I0(GND_net), .I1(n840_adj_1969[4]), 
            .I2(n331_adj_1114), .I3(n16381), .O(n839_adj_1968[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_7 (.CI(n16381), .I0(n840_adj_1969[4]), .I1(n331_adj_1114), 
            .CO(n16382));
    SB_LUT4 D_15__I_0_add_568_6_lut (.I0(GND_net), .I1(n840_adj_1969[3]), 
            .I2(n282_adj_1116), .I3(n16380), .O(n839_adj_1968[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_6 (.CI(n16380), .I0(n840_adj_1969[3]), .I1(n282_adj_1116), 
            .CO(n16381));
    SB_LUT4 D_15__I_0_add_568_5_lut (.I0(GND_net), .I1(n840_adj_1969[2]), 
            .I2(n233), .I3(n16379), .O(n839_adj_1968[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_5 (.CI(n16379), .I0(n840_adj_1969[2]), .I1(n233), 
            .CO(n16380));
    SB_LUT4 D_15__I_0_add_568_4_lut (.I0(GND_net), .I1(n840_adj_1969[1]), 
            .I2(n184_adj_1120), .I3(n16378), .O(n839_adj_1968[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_4 (.CI(n16378), .I0(n840_adj_1969[1]), .I1(n184_adj_1120), 
            .CO(n16379));
    SB_LUT4 D_15__I_0_add_568_3_lut (.I0(GND_net), .I1(n840_adj_1969[0]), 
            .I2(n135_adj_1123), .I3(n16377), .O(n839_adj_1968[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_3 (.CI(n16377), .I0(n840_adj_1969[0]), .I1(n135_adj_1123), 
            .CO(n16378));
    SB_LUT4 D_15__I_0_add_568_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n839_adj_1968[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_568_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16377));
    SB_LUT4 D_15__I_0_add_569_16_lut (.I0(GND_net), .I1(n841_adj_1970[13]), 
            .I2(n793_adj_1098), .I3(n16375), .O(n840_adj_1969[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_16 (.CI(n16375), .I0(n841_adj_1970[13]), 
            .I1(n793_adj_1098), .CO(n771_adj_1207));
    SB_LUT4 D_15__I_0_add_569_15_lut (.I0(GND_net), .I1(n841_adj_1970[12]), 
            .I2(n723_adj_1100), .I3(n16374), .O(n840_adj_1969[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_15 (.CI(n16374), .I0(n841_adj_1970[12]), 
            .I1(n723_adj_1100), .CO(n16375));
    SB_LUT4 D_15__I_0_add_569_14_lut (.I0(GND_net), .I1(n841_adj_1970[11]), 
            .I2(n674_adj_1101), .I3(n16373), .O(n840_adj_1969[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_14 (.CI(n16373), .I0(n841_adj_1970[11]), 
            .I1(n674_adj_1101), .CO(n16374));
    SB_LUT4 D_15__I_0_add_569_13_lut (.I0(GND_net), .I1(n841_adj_1970[10]), 
            .I2(n625_adj_1102), .I3(n16372), .O(n840_adj_1969[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_13 (.CI(n16372), .I0(n841_adj_1970[10]), 
            .I1(n625_adj_1102), .CO(n16373));
    SB_LUT4 D_15__I_0_add_569_12_lut (.I0(GND_net), .I1(n841_adj_1970[9]), 
            .I2(n576_adj_1104), .I3(n16371), .O(n840_adj_1969[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_12 (.CI(n16371), .I0(n841_adj_1970[9]), .I1(n576_adj_1104), 
            .CO(n16372));
    SB_LUT4 D_15__I_0_add_569_11_lut (.I0(GND_net), .I1(n841_adj_1970[8]), 
            .I2(n527_adj_1106), .I3(n16370), .O(n840_adj_1969[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_11 (.CI(n16370), .I0(n841_adj_1970[8]), .I1(n527_adj_1106), 
            .CO(n16371));
    SB_LUT4 D_15__I_0_add_569_10_lut (.I0(GND_net), .I1(n841_adj_1970[7]), 
            .I2(n478_adj_1108), .I3(n16369), .O(n840_adj_1969[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_10 (.CI(n16369), .I0(n841_adj_1970[7]), .I1(n478_adj_1108), 
            .CO(n16370));
    SB_CARRY Q_15__I_0_11_add_565_3 (.CI(n16631), .I0(n837_adj_1955[0]), 
            .I1(n135_c), .CO(n16632));
    SB_LUT4 D_15__I_0_add_569_9_lut (.I0(GND_net), .I1(n841_adj_1970[6]), 
            .I2(n429_adj_1110), .I3(n16368), .O(n840_adj_1969[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_9 (.CI(n16368), .I0(n841_adj_1970[6]), .I1(n429_adj_1110), 
            .CO(n16369));
    SB_LUT4 D_15__I_0_add_569_8_lut (.I0(GND_net), .I1(n841_adj_1970[5]), 
            .I2(n380_adj_1112), .I3(n16367), .O(n840_adj_1969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_9_lut (.I0(GND_net), .I1(n843_adj_1956[6]), 
            .I2(n423), .I3(n16741), .O(n842_adj_1954[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_8 (.CI(n16367), .I0(n841_adj_1970[5]), .I1(n380_adj_1112), 
            .CO(n16368));
    SB_LUT4 D_15__I_0_add_569_7_lut (.I0(GND_net), .I1(n841_adj_1970[4]), 
            .I2(n331_adj_1114), .I3(n16366), .O(n840_adj_1969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_7 (.CI(n16366), .I0(n841_adj_1970[4]), .I1(n331_adj_1114), 
            .CO(n16367));
    SB_LUT4 D_15__I_0_add_569_6_lut (.I0(GND_net), .I1(n841_adj_1970[3]), 
            .I2(n282_adj_1116), .I3(n16365), .O(n840_adj_1969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_6 (.CI(n16365), .I0(n841_adj_1970[3]), .I1(n282_adj_1116), 
            .CO(n16366));
    SB_LUT4 D_15__I_0_add_569_5_lut (.I0(GND_net), .I1(n841_adj_1970[2]), 
            .I2(n233), .I3(n16364), .O(n840_adj_1969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_5 (.CI(n16364), .I0(n841_adj_1970[2]), .I1(n233), 
            .CO(n16365));
    SB_CARRY D_15__I_0_10_add_571_9 (.CI(n16741), .I0(n843_adj_1956[6]), 
            .I1(n423), .CO(n16742));
    SB_LUT4 D_15__I_0_add_569_4_lut (.I0(GND_net), .I1(n841_adj_1970[1]), 
            .I2(n184_adj_1120), .I3(n16363), .O(n840_adj_1969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_4 (.CI(n16363), .I0(n841_adj_1970[1]), .I1(n184_adj_1120), 
            .CO(n16364));
    SB_LUT4 D_15__I_0_add_569_3_lut (.I0(GND_net), .I1(n841_adj_1970[0]), 
            .I2(n135_adj_1123), .I3(n16362), .O(n840_adj_1969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_3 (.CI(n16362), .I0(n841_adj_1970[0]), .I1(n135_adj_1123), 
            .CO(n16363));
    SB_LUT4 D_15__I_0_add_569_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n840_adj_1969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_569_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16362));
    SB_LUT4 D_15__I_0_add_570_16_lut (.I0(GND_net), .I1(n842_adj_1971[13]), 
            .I2(n793_adj_1098), .I3(n16360), .O(n841_adj_1970[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_16 (.CI(n16360), .I0(n842_adj_1971[13]), 
            .I1(n793_adj_1098), .CO(n775_adj_1224));
    SB_LUT4 D_15__I_0_add_570_15_lut (.I0(GND_net), .I1(n842_adj_1971[12]), 
            .I2(n723_adj_1100), .I3(n16359), .O(n841_adj_1970[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_15 (.CI(n16359), .I0(n842_adj_1971[12]), 
            .I1(n723_adj_1100), .CO(n16360));
    SB_LUT4 D_15__I_0_add_570_14_lut (.I0(GND_net), .I1(n842_adj_1971[11]), 
            .I2(n674_adj_1101), .I3(n16358), .O(n841_adj_1970[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_8_lut (.I0(GND_net), .I1(n843_adj_1956[5]), 
            .I2(n374), .I3(n16740), .O(n842_adj_1954[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_8 (.CI(n16740), .I0(n843_adj_1956[5]), 
            .I1(n374), .CO(n16741));
    SB_CARRY D_15__I_0_add_570_14 (.CI(n16358), .I0(n842_adj_1971[11]), 
            .I1(n674_adj_1101), .CO(n16359));
    SB_LUT4 D_15__I_0_add_570_13_lut (.I0(GND_net), .I1(n842_adj_1971[10]), 
            .I2(n625_adj_1102), .I3(n16357), .O(n841_adj_1970[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_13 (.CI(n16357), .I0(n842_adj_1971[10]), 
            .I1(n625_adj_1102), .CO(n16358));
    SB_LUT4 D_15__I_0_add_570_12_lut (.I0(GND_net), .I1(n842_adj_1971[9]), 
            .I2(n576_adj_1104), .I3(n16356), .O(n841_adj_1970[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_12 (.CI(n16356), .I0(n842_adj_1971[9]), .I1(n576_adj_1104), 
            .CO(n16357));
    SB_LUT4 D_15__I_0_add_570_11_lut (.I0(GND_net), .I1(n842_adj_1971[8]), 
            .I2(n527_adj_1106), .I3(n16355), .O(n841_adj_1970[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_11 (.CI(n16355), .I0(n842_adj_1971[8]), .I1(n527_adj_1106), 
            .CO(n16356));
    SB_LUT4 D_15__I_0_add_570_10_lut (.I0(GND_net), .I1(n842_adj_1971[7]), 
            .I2(n478_adj_1108), .I3(n16354), .O(n841_adj_1970[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_10 (.CI(n16354), .I0(n842_adj_1971[7]), .I1(n478_adj_1108), 
            .CO(n16355));
    SB_LUT4 D_15__I_0_add_570_9_lut (.I0(GND_net), .I1(n842_adj_1971[6]), 
            .I2(n429_adj_1110), .I3(n16353), .O(n841_adj_1970[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_9 (.CI(n16353), .I0(n842_adj_1971[6]), .I1(n429_adj_1110), 
            .CO(n16354));
    SB_LUT4 D_15__I_0_add_570_8_lut (.I0(GND_net), .I1(n842_adj_1971[5]), 
            .I2(n380_adj_1112), .I3(n16352), .O(n841_adj_1970[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_8 (.CI(n16352), .I0(n842_adj_1971[5]), .I1(n380_adj_1112), 
            .CO(n16353));
    SB_LUT4 D_15__I_0_add_570_7_lut (.I0(GND_net), .I1(n842_adj_1971[4]), 
            .I2(n331_adj_1114), .I3(n16351), .O(n841_adj_1970[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_7 (.CI(n16351), .I0(n842_adj_1971[4]), .I1(n331_adj_1114), 
            .CO(n16352));
    SB_LUT4 D_15__I_0_add_570_6_lut (.I0(GND_net), .I1(n842_adj_1971[3]), 
            .I2(n282_adj_1116), .I3(n16350), .O(n841_adj_1970[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_6 (.CI(n16350), .I0(n842_adj_1971[3]), .I1(n282_adj_1116), 
            .CO(n16351));
    SB_LUT4 D_15__I_0_add_570_5_lut (.I0(GND_net), .I1(n842_adj_1971[2]), 
            .I2(n233), .I3(n16349), .O(n841_adj_1970[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_5 (.CI(n16349), .I0(n842_adj_1971[2]), .I1(n233), 
            .CO(n16350));
    SB_LUT4 D_15__I_0_add_570_4_lut (.I0(GND_net), .I1(n842_adj_1971[1]), 
            .I2(n184_adj_1120), .I3(n16348), .O(n841_adj_1970[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_4 (.CI(n16348), .I0(n842_adj_1971[1]), .I1(n184_adj_1120), 
            .CO(n16349));
    SB_LUT4 D_15__I_0_add_570_3_lut (.I0(GND_net), .I1(n842_adj_1971[0]), 
            .I2(n135_adj_1123), .I3(n16347), .O(n841_adj_1970[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_3 (.CI(n16347), .I0(n842_adj_1971[0]), .I1(n135_adj_1123), 
            .CO(n16348));
    SB_LUT4 D_15__I_0_add_570_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n841_adj_1970[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_570_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16347));
    SB_LUT4 D_15__I_0_add_571_16_lut (.I0(GND_net), .I1(n843_adj_1972[13]), 
            .I2(n793_adj_1098), .I3(n16345), .O(n842_adj_1971[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_16 (.CI(n16345), .I0(n843_adj_1972[13]), 
            .I1(n793_adj_1098), .CO(n779_adj_1241));
    SB_LUT4 D_15__I_0_add_571_15_lut (.I0(GND_net), .I1(n843_adj_1972[12]), 
            .I2(n723_adj_1100), .I3(n16344), .O(n842_adj_1971[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_15 (.CI(n16344), .I0(n843_adj_1972[12]), 
            .I1(n723_adj_1100), .CO(n16345));
    SB_LUT4 D_15__I_0_add_571_14_lut (.I0(GND_net), .I1(n843_adj_1972[11]), 
            .I2(n674_adj_1101), .I3(n16343), .O(n842_adj_1971[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_14 (.CI(n16343), .I0(n843_adj_1972[11]), 
            .I1(n674_adj_1101), .CO(n16344));
    SB_LUT4 D_15__I_0_add_571_13_lut (.I0(GND_net), .I1(n843_adj_1972[10]), 
            .I2(n625_adj_1102), .I3(n16342), .O(n842_adj_1971[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_13 (.CI(n16342), .I0(n843_adj_1972[10]), 
            .I1(n625_adj_1102), .CO(n16343));
    SB_LUT4 D_15__I_0_add_571_12_lut (.I0(GND_net), .I1(n843_adj_1972[9]), 
            .I2(n576_adj_1104), .I3(n16341), .O(n842_adj_1971[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_12 (.CI(n16341), .I0(n843_adj_1972[9]), .I1(n576_adj_1104), 
            .CO(n16342));
    SB_LUT4 D_15__I_0_add_571_11_lut (.I0(GND_net), .I1(n843_adj_1972[8]), 
            .I2(n527_adj_1106), .I3(n16340), .O(n842_adj_1971[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_11 (.CI(n16340), .I0(n843_adj_1972[8]), .I1(n527_adj_1106), 
            .CO(n16341));
    SB_LUT4 D_15__I_0_add_571_10_lut (.I0(GND_net), .I1(n843_adj_1972[7]), 
            .I2(n478_adj_1108), .I3(n16339), .O(n842_adj_1971[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_10 (.CI(n16339), .I0(n843_adj_1972[7]), .I1(n478_adj_1108), 
            .CO(n16340));
    SB_LUT4 D_15__I_0_add_571_9_lut (.I0(GND_net), .I1(n843_adj_1972[6]), 
            .I2(n429_adj_1110), .I3(n16338), .O(n842_adj_1971[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_9 (.CI(n16338), .I0(n843_adj_1972[6]), .I1(n429_adj_1110), 
            .CO(n16339));
    SB_LUT4 D_15__I_0_add_571_8_lut (.I0(GND_net), .I1(n843_adj_1972[5]), 
            .I2(n380_adj_1112), .I3(n16337), .O(n842_adj_1971[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_8 (.CI(n16337), .I0(n843_adj_1972[5]), .I1(n380_adj_1112), 
            .CO(n16338));
    SB_LUT4 D_15__I_0_add_571_7_lut (.I0(GND_net), .I1(n843_adj_1972[4]), 
            .I2(n331_adj_1114), .I3(n16336), .O(n842_adj_1971[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_7 (.CI(n16336), .I0(n843_adj_1972[4]), .I1(n331_adj_1114), 
            .CO(n16337));
    SB_LUT4 D_15__I_0_add_571_6_lut (.I0(GND_net), .I1(n843_adj_1972[3]), 
            .I2(n282_adj_1116), .I3(n16335), .O(n842_adj_1971[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_6 (.CI(n16335), .I0(n843_adj_1972[3]), .I1(n282_adj_1116), 
            .CO(n16336));
    SB_LUT4 D_15__I_0_add_571_5_lut (.I0(GND_net), .I1(n843_adj_1972[2]), 
            .I2(n233), .I3(n16334), .O(n842_adj_1971[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_5 (.CI(n16334), .I0(n843_adj_1972[2]), .I1(n233), 
            .CO(n16335));
    SB_LUT4 D_15__I_0_add_571_4_lut (.I0(GND_net), .I1(n843_adj_1972[1]), 
            .I2(n184_adj_1120), .I3(n16333), .O(n842_adj_1971[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_4 (.CI(n16333), .I0(n843_adj_1972[1]), .I1(n184_adj_1120), 
            .CO(n16334));
    SB_LUT4 D_15__I_0_add_571_3_lut (.I0(GND_net), .I1(n843_adj_1972[0]), 
            .I2(n135_adj_1123), .I3(n16332), .O(n842_adj_1971[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_3 (.CI(n16332), .I0(n843_adj_1972[0]), .I1(n135_adj_1123), 
            .CO(n16333));
    SB_LUT4 D_15__I_0_add_571_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n842_adj_1971[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_571_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16332));
    SB_LUT4 D_15__I_0_add_572_16_lut (.I0(GND_net), .I1(n844_adj_1973[13]), 
            .I2(n793_adj_1098), .I3(n16330), .O(n843_adj_1972[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_16 (.CI(n16330), .I0(n844_adj_1973[13]), 
            .I1(n793_adj_1098), .CO(n783_adj_1257));
    SB_LUT4 D_15__I_0_add_572_15_lut (.I0(GND_net), .I1(n844_adj_1973[12]), 
            .I2(n723_adj_1100), .I3(n16329), .O(n843_adj_1972[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_15 (.CI(n16329), .I0(n844_adj_1973[12]), 
            .I1(n723_adj_1100), .CO(n16330));
    SB_LUT4 D_15__I_0_add_572_14_lut (.I0(GND_net), .I1(n844_adj_1973[11]), 
            .I2(n674_adj_1101), .I3(n16328), .O(n843_adj_1972[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_14 (.CI(n16328), .I0(n844_adj_1973[11]), 
            .I1(n674_adj_1101), .CO(n16329));
    SB_LUT4 D_15__I_0_add_572_13_lut (.I0(GND_net), .I1(n844_adj_1973[10]), 
            .I2(n625_adj_1102), .I3(n16327), .O(n843_adj_1972[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_13 (.CI(n16327), .I0(n844_adj_1973[10]), 
            .I1(n625_adj_1102), .CO(n16328));
    SB_LUT4 D_15__I_0_add_572_12_lut (.I0(GND_net), .I1(n844_adj_1973[9]), 
            .I2(n576_adj_1104), .I3(n16326), .O(n843_adj_1972[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_12 (.CI(n16326), .I0(n844_adj_1973[9]), .I1(n576_adj_1104), 
            .CO(n16327));
    SB_LUT4 D_15__I_0_add_572_11_lut (.I0(GND_net), .I1(n844_adj_1973[8]), 
            .I2(n527_adj_1106), .I3(n16325), .O(n843_adj_1972[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_11 (.CI(n16325), .I0(n844_adj_1973[8]), .I1(n527_adj_1106), 
            .CO(n16326));
    SB_LUT4 D_15__I_0_add_572_10_lut (.I0(GND_net), .I1(n844_adj_1973[7]), 
            .I2(n478_adj_1108), .I3(n16324), .O(n843_adj_1972[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_10 (.CI(n16324), .I0(n844_adj_1973[7]), .I1(n478_adj_1108), 
            .CO(n16325));
    SB_LUT4 D_15__I_0_add_572_9_lut (.I0(GND_net), .I1(n844_adj_1973[6]), 
            .I2(n429_adj_1110), .I3(n16323), .O(n843_adj_1972[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_9 (.CI(n16323), .I0(n844_adj_1973[6]), .I1(n429_adj_1110), 
            .CO(n16324));
    SB_LUT4 D_15__I_0_add_572_8_lut (.I0(GND_net), .I1(n844_adj_1973[5]), 
            .I2(n380_adj_1112), .I3(n16322), .O(n843_adj_1972[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_8 (.CI(n16322), .I0(n844_adj_1973[5]), .I1(n380_adj_1112), 
            .CO(n16323));
    SB_LUT4 D_15__I_0_add_572_7_lut (.I0(GND_net), .I1(n844_adj_1973[4]), 
            .I2(n331_adj_1114), .I3(n16321), .O(n843_adj_1972[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_7 (.CI(n16321), .I0(n844_adj_1973[4]), .I1(n331_adj_1114), 
            .CO(n16322));
    SB_LUT4 D_15__I_0_add_572_6_lut (.I0(GND_net), .I1(n844_adj_1973[3]), 
            .I2(n282_adj_1116), .I3(n16320), .O(n843_adj_1972[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_6 (.CI(n16320), .I0(n844_adj_1973[3]), .I1(n282_adj_1116), 
            .CO(n16321));
    SB_LUT4 D_15__I_0_add_572_5_lut (.I0(GND_net), .I1(n844_adj_1973[2]), 
            .I2(n233), .I3(n16319), .O(n843_adj_1972[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_5 (.CI(n16319), .I0(n844_adj_1973[2]), .I1(n233), 
            .CO(n16320));
    SB_LUT4 D_15__I_0_add_572_4_lut (.I0(GND_net), .I1(n844_adj_1973[1]), 
            .I2(n184_adj_1120), .I3(n16318), .O(n843_adj_1972[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_4 (.CI(n16318), .I0(n844_adj_1973[1]), .I1(n184_adj_1120), 
            .CO(n16319));
    SB_LUT4 D_15__I_0_add_572_3_lut (.I0(GND_net), .I1(n844_adj_1973[0]), 
            .I2(n135_adj_1123), .I3(n16317), .O(n843_adj_1972[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_3 (.CI(n16317), .I0(n844_adj_1973[0]), .I1(n135_adj_1123), 
            .CO(n16318));
    SB_LUT4 D_15__I_0_add_572_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n843_adj_1972[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_572_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16317));
    SB_LUT4 D_15__I_0_add_573_16_lut (.I0(GND_net), .I1(n845_adj_1974[13]), 
            .I2(n793_adj_1098), .I3(n16315), .O(n844_adj_1973[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_16 (.CI(n16315), .I0(n845_adj_1974[13]), 
            .I1(n793_adj_1098), .CO(n787_adj_1273));
    SB_LUT4 D_15__I_0_add_573_15_lut (.I0(GND_net), .I1(n845_adj_1974[12]), 
            .I2(n723_adj_1100), .I3(n16314), .O(n844_adj_1973[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_15 (.CI(n16314), .I0(n845_adj_1974[12]), 
            .I1(n723_adj_1100), .CO(n16315));
    SB_LUT4 D_15__I_0_add_573_14_lut (.I0(GND_net), .I1(n845_adj_1974[11]), 
            .I2(n674_adj_1101), .I3(n16313), .O(n844_adj_1973[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_14 (.CI(n16313), .I0(n845_adj_1974[11]), 
            .I1(n674_adj_1101), .CO(n16314));
    SB_LUT4 D_15__I_0_add_573_13_lut (.I0(GND_net), .I1(n845_adj_1974[10]), 
            .I2(n625_adj_1102), .I3(n16312), .O(n844_adj_1973[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_13 (.CI(n16312), .I0(n845_adj_1974[10]), 
            .I1(n625_adj_1102), .CO(n16313));
    SB_LUT4 D_15__I_0_add_573_12_lut (.I0(GND_net), .I1(n845_adj_1974[9]), 
            .I2(n576_adj_1104), .I3(n16311), .O(n844_adj_1973[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_12 (.CI(n16311), .I0(n845_adj_1974[9]), .I1(n576_adj_1104), 
            .CO(n16312));
    SB_LUT4 D_15__I_0_add_573_11_lut (.I0(GND_net), .I1(n845_adj_1974[8]), 
            .I2(n527_adj_1106), .I3(n16310), .O(n844_adj_1973[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_11 (.CI(n16310), .I0(n845_adj_1974[8]), .I1(n527_adj_1106), 
            .CO(n16311));
    SB_LUT4 D_15__I_0_add_573_10_lut (.I0(GND_net), .I1(n845_adj_1974[7]), 
            .I2(n478_adj_1108), .I3(n16309), .O(n844_adj_1973[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_10 (.CI(n16309), .I0(n845_adj_1974[7]), .I1(n478_adj_1108), 
            .CO(n16310));
    SB_LUT4 D_15__I_0_add_573_9_lut (.I0(GND_net), .I1(n845_adj_1974[6]), 
            .I2(n429_adj_1110), .I3(n16308), .O(n844_adj_1973[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_9 (.CI(n16308), .I0(n845_adj_1974[6]), .I1(n429_adj_1110), 
            .CO(n16309));
    SB_LUT4 D_15__I_0_add_573_8_lut (.I0(GND_net), .I1(n845_adj_1974[5]), 
            .I2(n380_adj_1112), .I3(n16307), .O(n844_adj_1973[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_8 (.CI(n16307), .I0(n845_adj_1974[5]), .I1(n380_adj_1112), 
            .CO(n16308));
    SB_LUT4 D_15__I_0_add_573_7_lut (.I0(GND_net), .I1(n845_adj_1974[4]), 
            .I2(n331_adj_1114), .I3(n16306), .O(n844_adj_1973[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_7 (.CI(n16306), .I0(n845_adj_1974[4]), .I1(n331_adj_1114), 
            .CO(n16307));
    SB_LUT4 D_15__I_0_add_573_6_lut (.I0(GND_net), .I1(n845_adj_1974[3]), 
            .I2(n282_adj_1116), .I3(n16305), .O(n844_adj_1973[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_6 (.CI(n16305), .I0(n845_adj_1974[3]), .I1(n282_adj_1116), 
            .CO(n16306));
    SB_LUT4 D_15__I_0_add_573_5_lut (.I0(GND_net), .I1(n845_adj_1974[2]), 
            .I2(n233), .I3(n16304), .O(n844_adj_1973[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_5 (.CI(n16304), .I0(n845_adj_1974[2]), .I1(n233), 
            .CO(n16305));
    SB_LUT4 D_15__I_0_add_573_4_lut (.I0(GND_net), .I1(n845_adj_1974[1]), 
            .I2(n184_adj_1120), .I3(n16303), .O(n844_adj_1973[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_4 (.CI(n16303), .I0(n845_adj_1974[1]), .I1(n184_adj_1120), 
            .CO(n16304));
    SB_LUT4 D_15__I_0_add_573_3_lut (.I0(GND_net), .I1(n845_adj_1974[0]), 
            .I2(n135_adj_1123), .I3(n16302), .O(n844_adj_1973[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_3 (.CI(n16302), .I0(n845_adj_1974[0]), .I1(n135_adj_1123), 
            .CO(n16303));
    SB_LUT4 D_15__I_0_add_573_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n844_adj_1973[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_573_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16302));
    SB_LUT4 D_15__I_0_add_574_16_lut (.I0(GND_net), .I1(n846_adj_1975[13]), 
            .I2(n793_adj_1098), .I3(n16300), .O(n845_adj_1974[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_16 (.CI(n16300), .I0(n846_adj_1975[13]), 
            .I1(n793_adj_1098), .CO(n791_adj_1289));
    SB_LUT4 D_15__I_0_add_574_15_lut (.I0(GND_net), .I1(n846_adj_1975[12]), 
            .I2(n723_adj_1100), .I3(n16299), .O(n845_adj_1974[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_15 (.CI(n16299), .I0(n846_adj_1975[12]), 
            .I1(n723_adj_1100), .CO(n16300));
    SB_LUT4 D_15__I_0_add_574_14_lut (.I0(GND_net), .I1(n846_adj_1975[11]), 
            .I2(n674_adj_1101), .I3(n16298), .O(n845_adj_1974[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_565_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n836[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_7_lut (.I0(GND_net), .I1(n843_adj_1956[4]), 
            .I2(n325), .I3(n16739), .O(n842_adj_1954[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_14 (.CI(n16298), .I0(n846_adj_1975[11]), 
            .I1(n674_adj_1101), .CO(n16299));
    SB_LUT4 D_15__I_0_add_574_13_lut (.I0(GND_net), .I1(n846_adj_1975[10]), 
            .I2(n625_adj_1102), .I3(n16297), .O(n845_adj_1974[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_13 (.CI(n16297), .I0(n846_adj_1975[10]), 
            .I1(n625_adj_1102), .CO(n16298));
    SB_LUT4 D_15__I_0_add_574_12_lut (.I0(GND_net), .I1(n846_adj_1975[9]), 
            .I2(n576_adj_1104), .I3(n16296), .O(n845_adj_1974[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_12 (.CI(n16296), .I0(n846_adj_1975[9]), .I1(n576_adj_1104), 
            .CO(n16297));
    SB_LUT4 D_15__I_0_add_574_11_lut (.I0(GND_net), .I1(n846_adj_1975[8]), 
            .I2(n527_adj_1106), .I3(n16295), .O(n845_adj_1974[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_7 (.CI(n16739), .I0(n843_adj_1956[4]), 
            .I1(n325), .CO(n16740));
    SB_CARRY D_15__I_0_add_574_11 (.CI(n16295), .I0(n846_adj_1975[8]), .I1(n527_adj_1106), 
            .CO(n16296));
    SB_LUT4 D_15__I_0_add_574_10_lut (.I0(GND_net), .I1(n846_adj_1975[7]), 
            .I2(n478_adj_1108), .I3(n16294), .O(n845_adj_1974[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_10 (.CI(n16294), .I0(n846_adj_1975[7]), .I1(n478_adj_1108), 
            .CO(n16295));
    SB_LUT4 D_15__I_0_add_574_9_lut (.I0(GND_net), .I1(n846_adj_1975[6]), 
            .I2(n429_adj_1110), .I3(n16293), .O(n845_adj_1974[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_9 (.CI(n16293), .I0(n846_adj_1975[6]), .I1(n429_adj_1110), 
            .CO(n16294));
    SB_LUT4 D_15__I_0_add_574_8_lut (.I0(GND_net), .I1(n846_adj_1975[5]), 
            .I2(n380_adj_1112), .I3(n16292), .O(n845_adj_1974[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_8 (.CI(n16292), .I0(n846_adj_1975[5]), .I1(n380_adj_1112), 
            .CO(n16293));
    SB_LUT4 D_15__I_0_add_574_7_lut (.I0(GND_net), .I1(n846_adj_1975[4]), 
            .I2(n331_adj_1114), .I3(n16291), .O(n845_adj_1974[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_7 (.CI(n16291), .I0(n846_adj_1975[4]), .I1(n331_adj_1114), 
            .CO(n16292));
    SB_LUT4 D_15__I_0_add_574_6_lut (.I0(GND_net), .I1(n846_adj_1975[3]), 
            .I2(n282_adj_1116), .I3(n16290), .O(n845_adj_1974[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_6 (.CI(n16290), .I0(n846_adj_1975[3]), .I1(n282_adj_1116), 
            .CO(n16291));
    SB_LUT4 D_15__I_0_10_add_571_6_lut (.I0(GND_net), .I1(n843_adj_1956[3]), 
            .I2(n276), .I3(n16738), .O(n842_adj_1954[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_6 (.CI(n16738), .I0(n843_adj_1956[3]), 
            .I1(n276), .CO(n16739));
    SB_LUT4 D_15__I_0_add_574_5_lut (.I0(GND_net), .I1(n846_adj_1975[2]), 
            .I2(n233), .I3(n16289), .O(n845_adj_1974[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_5 (.CI(n16289), .I0(n846_adj_1975[2]), .I1(n233), 
            .CO(n16290));
    SB_LUT4 D_15__I_0_add_574_4_lut (.I0(GND_net), .I1(n846_adj_1975[1]), 
            .I2(n184_adj_1120), .I3(n16288), .O(n845_adj_1974[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_4 (.CI(n16288), .I0(n846_adj_1975[1]), .I1(n184_adj_1120), 
            .CO(n16289));
    SB_LUT4 D_15__I_0_add_574_3_lut (.I0(GND_net), .I1(n846_adj_1975[0]), 
            .I2(n135_adj_1123), .I3(n16287), .O(n845_adj_1974[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_3 (.CI(n16287), .I0(n846_adj_1975[0]), .I1(n135_adj_1123), 
            .CO(n16288));
    SB_LUT4 D_15__I_0_add_574_2_lut (.I0(GND_net), .I1(\Product3_mul_temp[2] ), 
            .I2(n86_adj_204), .I3(GND_net), .O(n845_adj_1974[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_574_2 (.CI(GND_net), .I0(\Product3_mul_temp[2] ), 
            .I1(n86_adj_204), .CO(n16287));
    SB_LUT4 D_15__I_0_10_add_571_5_lut (.I0(GND_net), .I1(n843_adj_1956[2]), 
            .I2(n227), .I3(n16737), .O(n842_adj_1954[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_add_575_16_lut (.I0(GND_net), .I1(n19585), .I2(n793_adj_1098), 
            .I3(n16286), .O(n846_adj_1975[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_568_14_lut (.I0(GND_net), .I1(n840[11]), .I2(n674), 
            .I3(n16597), .O(n839[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_12_lut (.I0(GND_net), .I1(n538), .I2(n582_c), 
            .I3(n16685), .O(n846[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_add_575_15_lut (.I0(GND_net), .I1(n685_adj_205), .I2(n723_adj_1100), 
            .I3(n16285), .O(n846_adj_1975[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_15 (.CI(n16285), .I0(n685_adj_205), .I1(n723_adj_1100), 
            .CO(n16286));
    SB_LUT4 D_15__I_0_add_575_14_lut (.I0(GND_net), .I1(n636_adj_1310), 
            .I2(n674_adj_1101), .I3(n16284), .O(n846_adj_1975[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_14 (.CI(n16284), .I0(n636_adj_1310), .I1(n674_adj_1101), 
            .CO(n16285));
    SB_LUT4 D_15__I_0_add_575_13_lut (.I0(GND_net), .I1(n587_adj_206), .I2(n625_adj_1102), 
            .I3(n16283), .O(n846_adj_1975[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_13 (.CI(n16283), .I0(n587_adj_206), .I1(n625_adj_1102), 
            .CO(n16284));
    SB_LUT4 D_15__I_0_add_575_12_lut (.I0(GND_net), .I1(n538_adj_1312), 
            .I2(n576_adj_1104), .I3(n16282), .O(n846_adj_1975[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_12 (.CI(n16282), .I0(n538_adj_1312), .I1(n576_adj_1104), 
            .CO(n16283));
    SB_LUT4 Q_15__I_0_i101_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n148));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_add_575_11_lut (.I0(GND_net), .I1(n489_adj_207), .I2(n527_adj_1106), 
            .I3(n16281), .O(n846_adj_1975[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i134_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n197_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_add_575_11 (.CI(n16281), .I0(n489_adj_207), .I1(n527_adj_1106), 
            .CO(n16282));
    SB_LUT4 D_15__I_0_add_575_10_lut (.I0(GND_net), .I1(n440_adj_1314), 
            .I2(n478_adj_1108), .I3(n16280), .O(n846_adj_1975[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_10 (.CI(n16280), .I0(n440_adj_1314), .I1(n478_adj_1108), 
            .CO(n16281));
    SB_LUT4 D_15__I_0_add_575_9_lut (.I0(GND_net), .I1(n391_adj_208), .I2(n429_adj_1110), 
            .I3(n16279), .O(n846_adj_1975[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_9 (.CI(n16279), .I0(n391_adj_208), .I1(n429_adj_1110), 
            .CO(n16280));
    SB_LUT4 D_15__I_0_add_575_8_lut (.I0(GND_net), .I1(n342_adj_209), .I2(n380_adj_1112), 
            .I3(n16278), .O(n846_adj_1975[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_5 (.CI(n16737), .I0(n843_adj_1956[2]), 
            .I1(n227), .CO(n16738));
    SB_CARRY D_15__I_0_add_575_8 (.CI(n16278), .I0(n342_adj_209), .I1(n380_adj_1112), 
            .CO(n16279));
    SB_LUT4 D_15__I_0_add_575_7_lut (.I0(GND_net), .I1(n293_adj_1317), .I2(n331_adj_1114), 
            .I3(n16277), .O(n846_adj_1975[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_7 (.CI(n16277), .I0(n293_adj_1317), .I1(n331_adj_1114), 
            .CO(n16278));
    SB_CARRY Q_15__I_0_11_add_565_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16631));
    SB_LUT4 D_15__I_0_10_add_571_4_lut (.I0(GND_net), .I1(n843_adj_1956[1]), 
            .I2(n178), .I3(n16736), .O(n842_adj_1954[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_add_575_6_lut (.I0(GND_net), .I1(n244), .I2(n282_adj_1116), 
            .I3(n16276), .O(n846_adj_1975[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_6 (.CI(n16276), .I0(n244), .I1(n282_adj_1116), 
            .CO(n16277));
    SB_CARRY D_15__I_0_10_add_571_4 (.CI(n16736), .I0(n843_adj_1956[1]), 
            .I1(n178), .CO(n16737));
    SB_LUT4 D_15__I_0_add_575_5_lut (.I0(GND_net), .I1(n195_adj_1320), .I2(n233), 
            .I3(n16275), .O(n846_adj_1975[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_5 (.CI(n16275), .I0(n195_adj_1320), .I1(n233), 
            .CO(n16276));
    SB_LUT4 D_15__I_0_add_575_4_lut (.I0(GND_net), .I1(n146_adj_1321), .I2(n184_adj_1120), 
            .I3(n16274), .O(n846_adj_1975[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_4 (.CI(n16274), .I0(n146_adj_1321), .I1(n184_adj_1120), 
            .CO(n16275));
    SB_LUT4 D_15__I_0_add_575_3_lut (.I0(GND_net), .I1(n97_adj_1322), .I2(n135_adj_1123), 
            .I3(n16273), .O(n846_adj_1975[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_3 (.CI(n16273), .I0(n97_adj_1322), .I1(n135_adj_1123), 
            .CO(n16274));
    SB_LUT4 Q_15__I_0_11_add_566_16_lut (.I0(GND_net), .I1(n838_adj_1953[13]), 
            .I2(n793), .I3(n16629), .O(n837_adj_1955[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_571_3_lut (.I0(GND_net), .I1(n843_adj_1956[0]), 
            .I2(n129), .I3(n16735), .O(n842_adj_1954[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_add_575_2_lut (.I0(GND_net), .I1(n48_adj_1326), .I2(n86_adj_204), 
            .I3(GND_net), .O(n846_adj_1975[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_add_575_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_add_575_2 (.CI(GND_net), .I0(n48_adj_1326), .I1(n86_adj_204), 
            .CO(n16273));
    SB_LUT4 add_1229_16_lut (.I0(GND_net), .I1(n846_adj_1958[14]), .I2(n791), 
            .I3(n16272), .O(Product2_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_571_3 (.CI(n16735), .I0(n843_adj_1956[0]), 
            .I1(n129), .CO(n16736));
    SB_LUT4 add_1229_15_lut (.I0(GND_net), .I1(n845_adj_1957[14]), .I2(n787), 
            .I3(n16271), .O(Product2_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_16 (.CI(n16629), .I0(n838_adj_1953[13]), 
            .I1(n793), .CO(n759_adj_1327));
    SB_LUT4 D_15__I_0_10_add_571_2_lut (.I0(GND_net), .I1(n35), .I2(n80), 
            .I3(GND_net), .O(n842_adj_1954[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i200_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n295));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_1229_15 (.CI(n16271), .I0(n845_adj_1957[14]), .I1(n787), 
            .CO(n16272));
    SB_LUT4 add_1229_14_lut (.I0(GND_net), .I1(n844[14]), .I2(n783), .I3(n16270), 
            .O(Product2_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_14 (.CI(n16270), .I0(n844[14]), .I1(n783), .CO(n16271));
    SB_CARRY D_15__I_0_10_add_571_2 (.CI(GND_net), .I0(n35), .I1(n80), 
            .CO(n16735));
    SB_CARRY D_15__I_0_10_add_575_12 (.CI(n16685), .I0(n538), .I1(n582_c), 
            .CO(n16686));
    SB_LUT4 add_1229_13_lut (.I0(GND_net), .I1(n843[14]), .I2(n779), .I3(n16269), 
            .O(Product2_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_13 (.CI(n16269), .I0(n843[14]), .I1(n779), .CO(n16270));
    SB_LUT4 D_15__I_0_10_add_572_16_lut (.I0(GND_net), .I1(n844_adj_1959[13]), 
            .I2(n781), .I3(n16733), .O(n843_adj_1956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1229_12_lut (.I0(GND_net), .I1(n842[14]), .I2(n775_adj_1064), 
            .I3(n16268), .O(Product2_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_12 (.CI(n16268), .I0(n842[14]), .I1(n775_adj_1064), 
            .CO(n16269));
    SB_LUT4 Q_15__I_0_i233_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i299_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i299_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i332_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n491_adj_1330));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i332_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_1229_11_lut (.I0(GND_net), .I1(n841_adj_1952[14]), .I2(n771_adj_1019), 
            .I3(n16267), .O(Product2_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_11 (.CI(n16267), .I0(n841_adj_1952[14]), .I1(n771_adj_1019), 
            .CO(n16268));
    SB_LUT4 add_1229_10_lut (.I0(GND_net), .I1(n840[14]), .I2(n767), .I3(n16266), 
            .O(Product2_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_16 (.CI(n16733), .I0(n844_adj_1959[13]), 
            .I1(n781), .CO(n783_adj_1090));
    SB_CARRY add_1229_10 (.CI(n16266), .I0(n840[14]), .I1(n767), .CO(n16267));
    SB_LUT4 add_1229_9_lut (.I0(GND_net), .I1(n839[14]), .I2(n763_adj_1331), 
            .I3(n16265), .O(Product2_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_9 (.CI(n16265), .I0(n839[14]), .I1(n763_adj_1331), 
            .CO(n16266));
    SB_LUT4 add_1229_8_lut (.I0(GND_net), .I1(n838_adj_1953[14]), .I2(n759_adj_1327), 
            .I3(n16264), .O(Product2_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i431_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n638));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i431_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i200_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n295_adj_1333));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_1229_8 (.CI(n16264), .I0(n838_adj_1953[14]), .I1(n759_adj_1327), 
            .CO(n16265));
    SB_LUT4 add_1229_7_lut (.I0(GND_net), .I1(n837_adj_1955[14]), .I2(n755), 
            .I3(n16263), .O(Product2_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_7 (.CI(n16263), .I0(n837_adj_1955[14]), .I1(n755), 
            .CO(n16264));
    SB_LUT4 add_1229_6_lut (.I0(GND_net), .I1(n836[14]), .I2(n751_adj_1334), 
            .I3(n16262), .O(Product2_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_572_15_lut (.I0(GND_net), .I1(n844_adj_1959[12]), 
            .I2(n720), .I3(n16732), .O(n843_adj_1956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_6 (.CI(n16262), .I0(n836[14]), .I1(n751_adj_1334), 
            .CO(n16263));
    SB_CARRY D_15__I_0_10_add_572_15 (.CI(n16732), .I0(n844_adj_1959[12]), 
            .I1(n720), .CO(n16733));
    SB_LUT4 add_1229_5_lut (.I0(GND_net), .I1(n835[14]), .I2(n747_adj_1337), 
            .I3(n16261), .O(Product2_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_14 (.CI(n16597), .I0(n840[11]), .I1(n674), 
            .CO(n16598));
    SB_LUT4 D_15__I_0_10_add_575_11_lut (.I0(GND_net), .I1(n489_adj_210), 
            .I2(n533), .I3(n16684), .O(n846[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_568_13_lut (.I0(GND_net), .I1(n840[10]), .I2(n625_c), 
            .I3(n16596), .O(n839[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_11 (.CI(n16684), .I0(n489_adj_210), .I1(n533), 
            .CO(n16685));
    SB_CARRY Q_15__I_0_11_add_568_13 (.CI(n16596), .I0(n840[10]), .I1(n625_c), 
            .CO(n16597));
    SB_LUT4 D_15__I_0_10_add_575_10_lut (.I0(GND_net), .I1(n440_adj_1341), 
            .I2(n484), .I3(n16683), .O(n846[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_5 (.CI(n16261), .I0(n835[14]), .I1(n747_adj_1337), 
            .CO(n16262));
    SB_LUT4 Q_15__I_0_11_add_570_13_lut (.I0(GND_net), .I1(n842[10]), .I2(n625_c), 
            .I3(n16566), .O(n841_adj_1952[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1229_4_lut (.I0(GND_net), .I1(n834_adj_1976[14]), .I2(n9636), 
            .I3(n16260), .O(Product2_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_10 (.CI(n16683), .I0(n440_adj_1341), .I1(n484), 
            .CO(n16684));
    SB_CARRY add_1229_4 (.CI(n16260), .I0(n834_adj_1976[14]), .I1(n9636), 
            .CO(n16261));
    SB_LUT4 D_15__I_0_10_add_572_14_lut (.I0(GND_net), .I1(n844_adj_1959[11]), 
            .I2(n671), .I3(n16731), .O(n843_adj_1956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_566_15_lut (.I0(GND_net), .I1(n838_adj_1953[12]), 
            .I2(n723), .I3(n16628), .O(n837_adj_1955[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_14 (.CI(n16731), .I0(n844_adj_1959[11]), 
            .I1(n671), .CO(n16732));
    SB_LUT4 D_15__I_0_10_add_572_13_lut (.I0(GND_net), .I1(n844_adj_1959[10]), 
            .I2(n622), .I3(n16730), .O(n843_adj_1956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1229_3_lut (.I0(GND_net), .I1(n833_adj_1977[14]), .I2(n9213), 
            .I3(n16259), .O(Product2_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_568_14_lut (.I0(GND_net), .I1(n840_adj_1950[11]), 
            .I2(n659), .I3(n16791), .O(n839_adj_1951[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_6 (.CI(n16798), .I0(n839_adj_1951[3]), 
            .I1(n264), .CO(n16799));
    SB_LUT4 D_15__I_0_10_add_567_5_lut (.I0(GND_net), .I1(n839_adj_1951[2]), 
            .I2(n215), .I3(n16797), .O(n838[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_563_2 (.CI(GND_net), .I0(n11), .I1(n56), 
            .CO(n16855));
    SB_LUT4 D_15__I_0_10_add_564_16_lut (.I0(GND_net), .I1(n836_adj_1960[13]), 
            .I2(n749), .I3(n16853), .O(n835_adj_1961[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_3 (.CI(n16259), .I0(n833_adj_1977[14]), .I1(n9213), 
            .CO(n16260));
    SB_LUT4 add_1229_2_lut (.I0(GND_net), .I1(\qVoltage[15] ), .I2(\Product_mul_temp[26] ), 
            .I3(n16258), .O(Product2_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1229_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_2 (.CI(n16258), .I0(\qVoltage[15] ), .I1(\Product_mul_temp[26] ), 
            .CO(n16259));
    SB_CARRY D_15__I_0_10_add_563_11 (.CI(n16863), .I0(n835_adj_1961[8]), 
            .I1(n497_adj_1351), .CO(n16864));
    SB_LUT4 D_15__I_0_10_add_562_3_lut (.I0(GND_net), .I1(n834[0]), .I2(n102), 
            .I3(n16870), .O(n833[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1229_1 (.CI(GND_net), .I0(n832_adj_1978[14]), .I1(n832_adj_1978[14]), 
            .CO(n16258));
    SB_CARRY D_15__I_0_10_add_562_14 (.CI(n16881), .I0(n834[11]), .I1(n641_adj_1353), 
            .CO(n16882));
    SB_LUT4 add_1228_16_lut (.I0(GND_net), .I1(n846_adj_1975[14]), .I2(n791_adj_1289), 
            .I3(n16257), .O(Product3_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1228_15_lut (.I0(GND_net), .I1(n845_adj_1974[14]), .I2(n787_adj_1273), 
            .I3(n16256), .O(Product3_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_15 (.CI(n16256), .I0(n845_adj_1974[14]), .I1(n787_adj_1273), 
            .CO(n16257));
    SB_LUT4 add_1228_14_lut (.I0(GND_net), .I1(n844_adj_1973[14]), .I2(n783_adj_1257), 
            .I3(n16255), .O(Product3_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_562_13_lut (.I0(GND_net), .I1(n834[10]), .I2(n592), 
            .I3(n16880), .O(n833[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_9 (.CI(n16891), .I0(n833[6]), .I1(n393), 
            .CO(n16892));
    SB_LUT4 Q_15__I_0_11_add_568_12_lut (.I0(GND_net), .I1(n840[9]), .I2(n576), 
            .I3(n16595), .O(n839[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_9_lut (.I0(GND_net), .I1(n391_adj_211), 
            .I2(n435), .I3(n16682), .O(n846[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_14 (.CI(n16255), .I0(n844_adj_1973[14]), .I1(n783_adj_1257), 
            .CO(n16256));
    SB_LUT4 add_1228_13_lut (.I0(GND_net), .I1(n843_adj_1972[14]), .I2(n779_adj_1241), 
            .I3(n16254), .O(Product3_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_13 (.CI(n16254), .I0(n843_adj_1972[14]), .I1(n779_adj_1241), 
            .CO(n16255));
    SB_LUT4 add_1228_12_lut (.I0(GND_net), .I1(n842_adj_1971[14]), .I2(n775_adj_1224), 
            .I3(n16253), .O(Product3_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_12 (.CI(n16253), .I0(n842_adj_1971[14]), .I1(n775_adj_1224), 
            .CO(n16254));
    SB_LUT4 add_1228_11_lut (.I0(GND_net), .I1(n841_adj_1970[14]), .I2(n771_adj_1207), 
            .I3(n16252), .O(Product3_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_11 (.CI(n16252), .I0(n841_adj_1970[14]), .I1(n771_adj_1207), 
            .CO(n16253));
    SB_LUT4 add_1228_10_lut (.I0(GND_net), .I1(n840_adj_1969[14]), .I2(n767_adj_1191), 
            .I3(n16251), .O(Product3_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_10 (.CI(n16251), .I0(n840_adj_1969[14]), .I1(n767_adj_1191), 
            .CO(n16252));
    SB_LUT4 add_1228_9_lut (.I0(GND_net), .I1(n839_adj_1968[14]), .I2(n763_adj_1175), 
            .I3(n16250), .O(Product3_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_12 (.CI(n16595), .I0(n840[9]), .I1(n576), 
            .CO(n16596));
    SB_LUT4 D_15__I_0_10_add_566_12_lut (.I0(GND_net), .I1(n838[9]), .I2(n555_c), 
            .I3(n16819), .O(n837[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_9 (.CI(n16682), .I0(n391_adj_211), .I1(n435), 
            .CO(n16683));
    SB_CARRY D_15__I_0_10_add_566_12 (.CI(n16819), .I0(n838[9]), .I1(n555_c), 
            .CO(n16820));
    SB_LUT4 D_15__I_0_10_add_565_4_lut (.I0(GND_net), .I1(n837[1]), .I2(n160_adj_1359), 
            .I3(n16826), .O(n836_adj_1960[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_10 (.CI(n16832), .I0(n837[7]), .I1(n454_adj_1361), 
            .CO(n16833));
    SB_CARRY D_15__I_0_10_add_565_15 (.CI(n16837), .I0(n837[12]), .I1(n699_adj_1363), 
            .CO(n16838));
    SB_LUT4 D_15__I_0_10_add_565_14_lut (.I0(GND_net), .I1(n837[11]), .I2(n650_adj_1366), 
            .I3(n16836), .O(n836_adj_1960[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_6 (.CI(n16843), .I0(n836_adj_1960[3]), 
            .I1(n255), .CO(n16844));
    SB_LUT4 D_15__I_0_10_add_566_11_lut (.I0(GND_net), .I1(n838[8]), .I2(n506_adj_1370), 
            .I3(n16818), .O(n837[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_3 (.CI(n16810), .I0(n838[0]), .I1(n114), 
            .CO(n16811));
    SB_CARRY D_15__I_0_10_add_567_5 (.CI(n16797), .I0(n839_adj_1951[2]), 
            .I1(n215), .CO(n16798));
    SB_CARRY add_1228_9 (.CI(n16250), .I0(n839_adj_1968[14]), .I1(n763_adj_1175), 
            .CO(n16251));
    SB_LUT4 Q_15__I_0_11_add_568_11_lut (.I0(GND_net), .I1(n840[8]), .I2(n527), 
            .I3(n16594), .O(n839[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1228_8_lut (.I0(GND_net), .I1(n838_adj_1967[14]), .I2(n759_adj_1158), 
            .I3(n16249), .O(Product3_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_8 (.CI(n16249), .I0(n838_adj_1967[14]), .I1(n759_adj_1158), 
            .CO(n16250));
    SB_LUT4 add_1228_7_lut (.I0(GND_net), .I1(n837_adj_1966[14]), .I2(n755_adj_1144), 
            .I3(n16248), .O(Product3_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_13 (.CI(n16730), .I0(n844_adj_1959[10]), 
            .I1(n622), .CO(n16731));
    SB_CARRY add_1228_7 (.CI(n16248), .I0(n837_adj_1966[14]), .I1(n755_adj_1144), 
            .CO(n16249));
    SB_CARRY D_15__I_0_10_add_564_16 (.CI(n16853), .I0(n836_adj_1960[13]), 
            .I1(n749), .CO(n751));
    SB_LUT4 add_1228_6_lut (.I0(GND_net), .I1(n836_adj_1965[14]), .I2(n751_adj_1127), 
            .I3(n16247), .O(Product3_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_4_lut (.I0(GND_net), .I1(n839_adj_1951[1]), 
            .I2(n166), .I3(n16796), .O(n838[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_572_12_lut (.I0(GND_net), .I1(n844_adj_1959[9]), 
            .I2(n573_c), .I3(n16729), .O(n843_adj_1956[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_6 (.CI(n16247), .I0(n836_adj_1965[14]), .I1(n751_adj_1127), 
            .CO(n16248));
    SB_LUT4 add_1228_5_lut (.I0(GND_net), .I1(n835_adj_1963[14]), .I2(n747_adj_1099), 
            .I3(n16246), .O(Product3_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_10_lut (.I0(GND_net), .I1(n835_adj_1961[7]), 
            .I2(n448_adj_1374), .I3(n16862), .O(n834[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_3 (.CI(n16870), .I0(n834[0]), .I1(n102), 
            .CO(n16871));
    SB_CARRY D_15__I_0_10_add_562_13 (.CI(n16880), .I0(n834[10]), .I1(n592), 
            .CO(n16881));
    SB_LUT4 D_15__I_0_10_add_562_12_lut (.I0(GND_net), .I1(n834[9]), .I2(n543_c), 
            .I3(n16879), .O(n833[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_8_lut (.I0(GND_net), .I1(n342_adj_212), 
            .I2(n386), .I3(n16681), .O(n846[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_8_lut (.I0(GND_net), .I1(n833[5]), .I2(n344_adj_1377), 
            .I3(n16890), .O(Product1_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_16_lut (.I0(GND_net), .I1(n833[13]), .I2(n737), 
            .I3(n16898), .O(n832[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_564_15_lut (.I0(GND_net), .I1(n836_adj_1960[12]), 
            .I2(n696_adj_1380), .I3(n16852), .O(n835_adj_1961[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_11 (.CI(n16594), .I0(n840[8]), .I1(n527), 
            .CO(n16595));
    SB_CARRY add_1228_5 (.CI(n16246), .I0(n835_adj_1963[14]), .I1(n747_adj_1099), 
            .CO(n16247));
    SB_LUT4 add_1228_4_lut (.I0(GND_net), .I1(n834_adj_1962[14]), .I2(n9531), 
            .I3(n16245), .O(Product3_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_4 (.CI(n16245), .I0(n834_adj_1962[14]), .I1(n9531), 
            .CO(n16246));
    SB_LUT4 add_1228_3_lut (.I0(GND_net), .I1(n833_adj_1964[14]), .I2(n9108), 
            .I3(n16244), .O(Product3_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_3 (.CI(n16244), .I0(n833_adj_1964[14]), .I1(n9108), 
            .CO(n16245));
    SB_LUT4 add_1228_2_lut (.I0(GND_net), .I1(\dVoltage[15] ), .I2(\Product_mul_temp[26] ), 
            .I3(n16243), .O(Product3_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1228_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_2 (.CI(n16243), .I0(\dVoltage[15] ), .I1(\Product_mul_temp[26] ), 
            .CO(n16244));
    SB_CARRY D_15__I_0_10_add_572_12 (.CI(n16729), .I0(n844_adj_1959[9]), 
            .I1(n573_c), .CO(n16730));
    SB_CARRY D_15__I_0_10_add_575_8 (.CI(n16681), .I0(n342_adj_212), .I1(n386), 
            .CO(n16682));
    SB_LUT4 Q_15__I_0_11_add_568_10_lut (.I0(GND_net), .I1(n840[7]), .I2(n478), 
            .I3(n16593), .O(n839[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_12_lut (.I0(GND_net), .I1(n839_adj_1951[9]), 
            .I2(n558_c), .I3(n16804), .O(n838[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_12 (.CI(n16804), .I0(n839_adj_1951[9]), 
            .I1(n558_c), .CO(n16805));
    SB_LUT4 D_15__I_0_10_add_566_2_lut (.I0(GND_net), .I1(n20), .I2(n65), 
            .I3(GND_net), .O(n837[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_11 (.CI(n16818), .I0(n838[8]), .I1(n506_adj_1370), 
            .CO(n16819));
    SB_CARRY D_15__I_0_10_add_565_4 (.CI(n16826), .I0(n837[1]), .I1(n160_adj_1359), 
            .CO(n16827));
    SB_LUT4 D_15__I_0_10_add_565_3_lut (.I0(GND_net), .I1(n837[0]), .I2(n111), 
            .I3(n16825), .O(n836_adj_1960[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_7_lut (.I0(GND_net), .I1(n293_adj_1386), 
            .I2(n337), .I3(n16680), .O(n846[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1228_1 (.CI(GND_net), .I0(n832_adj_1979[14]), .I1(n832_adj_1979[14]), 
            .CO(n16243));
    SB_LUT4 D_15__I_0_10_add_565_9_lut (.I0(GND_net), .I1(n837[6]), .I2(n405), 
            .I3(n16831), .O(n836_adj_1960[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_15 (.CI(n16628), .I0(n838_adj_1953[12]), 
            .I1(n723), .CO(n16629));
    SB_CARRY D_15__I_0_10_add_565_14 (.CI(n16836), .I0(n837[11]), .I1(n650_adj_1366), 
            .CO(n16837));
    SB_LUT4 D_15__I_0_10_add_564_5_lut (.I0(GND_net), .I1(n836_adj_1960[2]), 
            .I2(n206), .I3(n16842), .O(n835_adj_1961[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_add_561_16_lut (.I0(GND_net), .I1(n833_adj_1981[13]), 
            .I2(n737_adj_213), .I3(n16241), .O(n832_adj_1980[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_572_11_lut (.I0(GND_net), .I1(n844_adj_1959[8]), 
            .I2(n524), .I3(n16728), .O(n843_adj_1956[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_5 (.CI(n16842), .I0(n836_adj_1960[2]), 
            .I1(n206), .CO(n16843));
    SB_LUT4 Q_15__I_0_11_add_566_14_lut (.I0(GND_net), .I1(n838_adj_1953[11]), 
            .I2(n674), .I3(n16627), .O(n837_adj_1955[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_14 (.CI(n16627), .I0(n838_adj_1953[11]), 
            .I1(n674), .CO(n16628));
    SB_LUT4 Q_15__I_0_11_add_566_13_lut (.I0(GND_net), .I1(n838_adj_1953[10]), 
            .I2(n625_c), .I3(n16626), .O(n837_adj_1955[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_16 (.CI(n16241), .I0(n833_adj_1981[13]), 
            .I1(n737_adj_213), .CO(n739_adj_1396));
    SB_LUT4 D_15__I_0_10_add_564_10_lut (.I0(GND_net), .I1(n836_adj_1960[7]), 
            .I2(n451_adj_1397), .I3(n16847), .O(n835_adj_1961[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_2 (.CI(GND_net), .I0(n20), .I1(n65), 
            .CO(n16810));
    SB_LUT4 D_15__I_0_10_add_564_13_lut (.I0(GND_net), .I1(n836_adj_1960[10]), 
            .I2(n598), .I3(n16850), .O(n835_adj_1961[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_11 (.CI(n16728), .I0(n844_adj_1959[8]), 
            .I1(n524), .CO(n16729));
    SB_LUT4 Q_15__I_0_add_561_15_lut (.I0(GND_net), .I1(n833_adj_1981[12]), 
            .I2(n687), .I3(n16240), .O(Product4_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_15 (.CI(n16852), .I0(n836_adj_1960[12]), 
            .I1(n696_adj_1380), .CO(n16853));
    SB_CARRY D_15__I_0_10_add_563_10 (.CI(n16862), .I0(n835_adj_1961[7]), 
            .I1(n448_adj_1374), .CO(n16863));
    SB_LUT4 D_15__I_0_10_add_563_9_lut (.I0(GND_net), .I1(n835_adj_1961[6]), 
            .I2(n399), .I3(n16861), .O(n834[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_562_2_lut (.I0(GND_net), .I1(n8), .I2(n53), 
            .I3(GND_net), .O(n833[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_12 (.CI(n16879), .I0(n834[9]), .I1(n543_c), 
            .CO(n16880));
    SB_CARRY D_15__I_0_10_add_561_8 (.CI(n16890), .I0(n833[5]), .I1(n344_adj_1377), 
            .CO(n16891));
    SB_LUT4 D_15__I_0_10_add_561_7_lut (.I0(GND_net), .I1(n833[4]), .I2(n295_adj_1333), 
            .I3(n16889), .O(Product1_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_16 (.CI(n16898), .I0(n833[13]), .I1(n737), 
            .CO(n739));
    SB_LUT4 Q_15__I_0_i464_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n687));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i305_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_1397));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i305_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i354_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i354_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_add_561_15 (.CI(n16240), .I0(n833_adj_1981[12]), 
            .I1(n687), .CO(n16241));
    SB_LUT4 Q_15__I_0_add_561_14_lut (.I0(GND_net), .I1(n833_adj_1981[11]), 
            .I2(n638), .I3(n16239), .O(Product4_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_14 (.CI(n16239), .I0(n833_adj_1981[11]), 
            .I1(n638), .CO(n16240));
    SB_LUT4 Q_15__I_0_add_561_13_lut (.I0(GND_net), .I1(n833_adj_1981[10]), 
            .I2(n589), .I3(n16238), .O(Product4_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_13 (.CI(n16238), .I0(n833_adj_1981[10]), 
            .I1(n589), .CO(n16239));
    SB_LUT4 Q_15__I_0_add_561_12_lut (.I0(GND_net), .I1(n833_adj_1981[9]), 
            .I2(n540), .I3(n16237), .O(Product4_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_12 (.CI(n16237), .I0(n833_adj_1981[9]), .I1(n540), 
            .CO(n16238));
    SB_LUT4 Q_15__I_0_add_561_11_lut (.I0(GND_net), .I1(n833_adj_1981[8]), 
            .I2(n491_adj_1330), .I3(n16236), .O(Product4_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_11 (.CI(n16236), .I0(n833_adj_1981[8]), .I1(n491_adj_1330), 
            .CO(n16237));
    SB_LUT4 Q_15__I_0_add_561_10_lut (.I0(GND_net), .I1(n833_adj_1981[7]), 
            .I2(n442), .I3(n16235), .O(Product4_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_10 (.CI(n16235), .I0(n833_adj_1981[7]), .I1(n442), 
            .CO(n16236));
    SB_LUT4 Q_15__I_0_add_561_9_lut (.I0(GND_net), .I1(n833_adj_1981[6]), 
            .I2(n393_adj_214), .I3(n16234), .O(Product4_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_9 (.CI(n16234), .I0(n833_adj_1981[6]), .I1(n393_adj_214), 
            .CO(n16235));
    SB_LUT4 Q_15__I_0_add_561_8_lut (.I0(GND_net), .I1(n833_adj_1981[5]), 
            .I2(n344), .I3(n16233), .O(Product4_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_8 (.CI(n16233), .I0(n833_adj_1981[5]), .I1(n344), 
            .CO(n16234));
    SB_LUT4 Q_15__I_0_add_561_7_lut (.I0(GND_net), .I1(n833_adj_1981[4]), 
            .I2(n295), .I3(n16232), .O(Product4_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_7 (.CI(n16232), .I0(n833_adj_1981[4]), .I1(n295), 
            .CO(n16233));
    SB_LUT4 Q_15__I_0_add_561_6_lut (.I0(GND_net), .I1(n833_adj_1981[3]), 
            .I2(n246), .I3(n16231), .O(Product4_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_6 (.CI(n16231), .I0(n833_adj_1981[3]), .I1(n246), 
            .CO(n16232));
    SB_LUT4 Q_15__I_0_add_561_5_lut (.I0(GND_net), .I1(n833_adj_1981[2]), 
            .I2(n197_c), .I3(n16230), .O(Product4_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_5 (.CI(n16230), .I0(n833_adj_1981[2]), .I1(n197_c), 
            .CO(n16231));
    SB_LUT4 Q_15__I_0_add_561_4_lut (.I0(GND_net), .I1(n833_adj_1981[1]), 
            .I2(n148), .I3(n16229), .O(Product4_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_4 (.CI(n16229), .I0(n833_adj_1981[1]), .I1(n148), 
            .CO(n16230));
    SB_LUT4 Q_15__I_0_add_561_3_lut (.I0(GND_net), .I1(n833_adj_1981[0]), 
            .I2(n99), .I3(n16228), .O(Product4_mul_temp[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_561_3 (.CI(n16228), .I0(n833_adj_1981[0]), .I1(n99), 
            .CO(n16229));
    SB_CARRY Q_15__I_0_add_561_2 (.CI(GND_net), .I0(n19351), .I1(n50), 
            .CO(n16228));
    SB_LUT4 Q_15__I_0_add_562_16_lut (.I0(GND_net), .I1(n834_adj_1982[13]), 
            .I2(n741), .I3(n16226), .O(n833_adj_1981[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_16 (.CI(n16226), .I0(n834_adj_1982[13]), 
            .I1(n741), .CO(n743_adj_1411));
    SB_LUT4 Q_15__I_0_add_562_15_lut (.I0(GND_net), .I1(n834_adj_1982[12]), 
            .I2(n690), .I3(n16225), .O(n833_adj_1981[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_15 (.CI(n16225), .I0(n834_adj_1982[12]), 
            .I1(n690), .CO(n16226));
    SB_LUT4 Q_15__I_0_add_562_14_lut (.I0(GND_net), .I1(n834_adj_1982[11]), 
            .I2(n641), .I3(n16224), .O(n833_adj_1981[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_14 (.CI(n16224), .I0(n834_adj_1982[11]), 
            .I1(n641), .CO(n16225));
    SB_LUT4 Q_15__I_0_add_562_13_lut (.I0(GND_net), .I1(n834_adj_1982[10]), 
            .I2(n592_adj_215), .I3(n16223), .O(n833_adj_1981[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_13 (.CI(n16223), .I0(n834_adj_1982[10]), 
            .I1(n592_adj_215), .CO(n16224));
    SB_LUT4 Q_15__I_0_add_562_12_lut (.I0(GND_net), .I1(n834_adj_1982[9]), 
            .I2(n543), .I3(n16222), .O(n833_adj_1981[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_12 (.CI(n16222), .I0(n834_adj_1982[9]), .I1(n543), 
            .CO(n16223));
    SB_LUT4 Q_15__I_0_add_562_11_lut (.I0(GND_net), .I1(n834_adj_1982[8]), 
            .I2(n494), .I3(n16221), .O(n833_adj_1981[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_11 (.CI(n16221), .I0(n834_adj_1982[8]), .I1(n494), 
            .CO(n16222));
    SB_LUT4 Q_15__I_0_add_562_10_lut (.I0(GND_net), .I1(n834_adj_1982[7]), 
            .I2(n445), .I3(n16220), .O(n833_adj_1981[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_10 (.CI(n16220), .I0(n834_adj_1982[7]), .I1(n445), 
            .CO(n16221));
    SB_LUT4 Q_15__I_0_add_562_9_lut (.I0(GND_net), .I1(n834_adj_1982[6]), 
            .I2(n396), .I3(n16219), .O(n833_adj_1981[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_9 (.CI(n16219), .I0(n834_adj_1982[6]), .I1(n396), 
            .CO(n16220));
    SB_LUT4 Q_15__I_0_add_562_8_lut (.I0(GND_net), .I1(n834_adj_1982[5]), 
            .I2(n347), .I3(n16218), .O(n833_adj_1981[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_8 (.CI(n16218), .I0(n834_adj_1982[5]), .I1(n347), 
            .CO(n16219));
    SB_LUT4 Q_15__I_0_add_562_7_lut (.I0(GND_net), .I1(n834_adj_1982[4]), 
            .I2(n298), .I3(n16217), .O(n833_adj_1981[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_7 (.CI(n16217), .I0(n834_adj_1982[4]), .I1(n298), 
            .CO(n16218));
    SB_LUT4 Q_15__I_0_add_562_6_lut (.I0(GND_net), .I1(n834_adj_1982[3]), 
            .I2(n249), .I3(n16216), .O(n833_adj_1981[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_6 (.CI(n16216), .I0(n834_adj_1982[3]), .I1(n249), 
            .CO(n16217));
    SB_LUT4 Q_15__I_0_add_562_5_lut (.I0(GND_net), .I1(n834_adj_1982[2]), 
            .I2(n200_c), .I3(n16215), .O(n833_adj_1981[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_5 (.CI(n16215), .I0(n834_adj_1982[2]), .I1(n200_c), 
            .CO(n16216));
    SB_LUT4 Q_15__I_0_add_562_4_lut (.I0(GND_net), .I1(n834_adj_1982[1]), 
            .I2(n151), .I3(n16214), .O(n833_adj_1981[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_4 (.CI(n16214), .I0(n834_adj_1982[1]), .I1(n151), 
            .CO(n16215));
    SB_LUT4 Q_15__I_0_add_562_3_lut (.I0(GND_net), .I1(n834_adj_1982[0]), 
            .I2(n102_adj_216), .I3(n16213), .O(n833_adj_1981[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_3 (.CI(n16213), .I0(n834_adj_1982[0]), .I1(n102_adj_216), 
            .CO(n16214));
    SB_LUT4 Q_15__I_0_add_562_2_lut (.I0(GND_net), .I1(n8_adj_217), .I2(n53_adj_218), 
            .I3(GND_net), .O(n833_adj_1981[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_562_2 (.CI(GND_net), .I0(n8_adj_217), .I1(n53_adj_218), 
            .CO(n16213));
    SB_LUT4 Q_15__I_0_add_563_16_lut (.I0(GND_net), .I1(n835_adj_1983[13]), 
            .I2(n745), .I3(n16211), .O(n834_adj_1982[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_16 (.CI(n16211), .I0(n835_adj_1983[13]), 
            .I1(n745), .CO(n747_adj_1425));
    SB_LUT4 Q_15__I_0_add_563_15_lut (.I0(GND_net), .I1(n835_adj_1983[12]), 
            .I2(n693), .I3(n16210), .O(n834_adj_1982[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_15 (.CI(n16210), .I0(n835_adj_1983[12]), 
            .I1(n693), .CO(n16211));
    SB_LUT4 Q_15__I_0_add_563_14_lut (.I0(GND_net), .I1(n835_adj_1983[11]), 
            .I2(n644), .I3(n16209), .O(n834_adj_1982[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_14 (.CI(n16209), .I0(n835_adj_1983[11]), 
            .I1(n644), .CO(n16210));
    SB_LUT4 Q_15__I_0_add_563_13_lut (.I0(GND_net), .I1(n835_adj_1983[10]), 
            .I2(n595), .I3(n16208), .O(n834_adj_1982[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_13 (.CI(n16208), .I0(n835_adj_1983[10]), 
            .I1(n595), .CO(n16209));
    SB_LUT4 Q_15__I_0_add_563_12_lut (.I0(GND_net), .I1(n835_adj_1983[9]), 
            .I2(n546), .I3(n16207), .O(n834_adj_1982[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_12 (.CI(n16207), .I0(n835_adj_1983[9]), .I1(n546), 
            .CO(n16208));
    SB_LUT4 Q_15__I_0_add_563_11_lut (.I0(GND_net), .I1(n835_adj_1983[8]), 
            .I2(n497), .I3(n16206), .O(n834_adj_1982[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_11 (.CI(n16206), .I0(n835_adj_1983[8]), .I1(n497), 
            .CO(n16207));
    SB_LUT4 Q_15__I_0_add_563_10_lut (.I0(GND_net), .I1(n835_adj_1983[7]), 
            .I2(n448), .I3(n16205), .O(n834_adj_1982[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_10 (.CI(n16205), .I0(n835_adj_1983[7]), .I1(n448), 
            .CO(n16206));
    SB_LUT4 Q_15__I_0_add_563_9_lut (.I0(GND_net), .I1(n835_adj_1983[6]), 
            .I2(n399_adj_219), .I3(n16204), .O(n834_adj_1982[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_9 (.CI(n16204), .I0(n835_adj_1983[6]), .I1(n399_adj_219), 
            .CO(n16205));
    SB_LUT4 Q_15__I_0_add_563_8_lut (.I0(GND_net), .I1(n835_adj_1983[5]), 
            .I2(n350), .I3(n16203), .O(n834_adj_1982[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_8 (.CI(n16203), .I0(n835_adj_1983[5]), .I1(n350), 
            .CO(n16204));
    SB_LUT4 Q_15__I_0_add_563_7_lut (.I0(GND_net), .I1(n835_adj_1983[4]), 
            .I2(n301), .I3(n16202), .O(n834_adj_1982[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_7 (.CI(n16202), .I0(n835_adj_1983[4]), .I1(n301), 
            .CO(n16203));
    SB_LUT4 Q_15__I_0_add_563_6_lut (.I0(GND_net), .I1(n835_adj_1983[3]), 
            .I2(n252), .I3(n16201), .O(n834_adj_1982[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_6 (.CI(n16201), .I0(n835_adj_1983[3]), .I1(n252), 
            .CO(n16202));
    SB_LUT4 Q_15__I_0_add_563_5_lut (.I0(GND_net), .I1(n835_adj_1983[2]), 
            .I2(n203_c), .I3(n16200), .O(n834_adj_1982[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_5 (.CI(n16200), .I0(n835_adj_1983[2]), .I1(n203_c), 
            .CO(n16201));
    SB_LUT4 Q_15__I_0_add_563_4_lut (.I0(GND_net), .I1(n835_adj_1983[1]), 
            .I2(n154), .I3(n16199), .O(n834_adj_1982[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_4 (.CI(n16199), .I0(n835_adj_1983[1]), .I1(n154), 
            .CO(n16200));
    SB_LUT4 Q_15__I_0_add_563_3_lut (.I0(GND_net), .I1(n835_adj_1983[0]), 
            .I2(n105), .I3(n16198), .O(n834_adj_1982[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_3 (.CI(n16198), .I0(n835_adj_1983[0]), .I1(n105), 
            .CO(n16199));
    SB_LUT4 Q_15__I_0_add_563_2_lut (.I0(GND_net), .I1(n11_adj_220), .I2(n56_adj_221), 
            .I3(GND_net), .O(n834_adj_1982[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_563_2 (.CI(GND_net), .I0(n11_adj_220), .I1(n56_adj_221), 
            .CO(n16198));
    SB_LUT4 Q_15__I_0_add_564_16_lut (.I0(GND_net), .I1(n836_adj_1984[13]), 
            .I2(n749_adj_222), .I3(n16196), .O(n835_adj_1983[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_16 (.CI(n16196), .I0(n836_adj_1984[13]), 
            .I1(n749_adj_222), .CO(n751_adj_1446));
    SB_LUT4 Q_15__I_0_add_564_15_lut (.I0(GND_net), .I1(n836_adj_1984[12]), 
            .I2(n696), .I3(n16195), .O(n835_adj_1983[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_15 (.CI(n16195), .I0(n836_adj_1984[12]), 
            .I1(n696), .CO(n16196));
    SB_LUT4 Q_15__I_0_add_564_14_lut (.I0(GND_net), .I1(n836_adj_1984[11]), 
            .I2(n647), .I3(n16194), .O(n835_adj_1983[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_14 (.CI(n16194), .I0(n836_adj_1984[11]), 
            .I1(n647), .CO(n16195));
    SB_LUT4 Q_15__I_0_add_564_13_lut (.I0(GND_net), .I1(n836_adj_1984[10]), 
            .I2(n598_adj_223), .I3(n16193), .O(n835_adj_1983[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_13 (.CI(n16193), .I0(n836_adj_1984[10]), 
            .I1(n598_adj_223), .CO(n16194));
    SB_LUT4 Q_15__I_0_add_564_12_lut (.I0(GND_net), .I1(n836_adj_1984[9]), 
            .I2(n549), .I3(n16192), .O(n835_adj_1983[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_12 (.CI(n16192), .I0(n836_adj_1984[9]), .I1(n549), 
            .CO(n16193));
    SB_LUT4 Q_15__I_0_add_564_11_lut (.I0(GND_net), .I1(n836_adj_1984[8]), 
            .I2(n500), .I3(n16191), .O(n835_adj_1983[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_11 (.CI(n16191), .I0(n836_adj_1984[8]), .I1(n500), 
            .CO(n16192));
    SB_LUT4 Q_15__I_0_add_564_10_lut (.I0(GND_net), .I1(n836_adj_1984[7]), 
            .I2(n451), .I3(n16190), .O(n835_adj_1983[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_10 (.CI(n16190), .I0(n836_adj_1984[7]), .I1(n451), 
            .CO(n16191));
    SB_LUT4 Q_15__I_0_add_564_9_lut (.I0(GND_net), .I1(n836_adj_1984[6]), 
            .I2(n402), .I3(n16189), .O(n835_adj_1983[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_9 (.CI(n16189), .I0(n836_adj_1984[6]), .I1(n402), 
            .CO(n16190));
    SB_LUT4 Q_15__I_0_add_564_8_lut (.I0(GND_net), .I1(n836_adj_1984[5]), 
            .I2(n353), .I3(n16188), .O(n835_adj_1983[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_8 (.CI(n16188), .I0(n836_adj_1984[5]), .I1(n353), 
            .CO(n16189));
    SB_LUT4 Q_15__I_0_add_564_7_lut (.I0(GND_net), .I1(n836_adj_1984[4]), 
            .I2(n304_adj_1031), .I3(n16187), .O(n835_adj_1983[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_7 (.CI(n16187), .I0(n836_adj_1984[4]), .I1(n304_adj_1031), 
            .CO(n16188));
    SB_LUT4 Q_15__I_0_add_564_6_lut (.I0(GND_net), .I1(n836_adj_1984[3]), 
            .I2(n255_adj_224), .I3(n16186), .O(n835_adj_1983[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_6 (.CI(n16186), .I0(n836_adj_1984[3]), .I1(n255_adj_224), 
            .CO(n16187));
    SB_LUT4 Q_15__I_0_add_564_5_lut (.I0(GND_net), .I1(n836_adj_1984[2]), 
            .I2(n206_c), .I3(n16185), .O(n835_adj_1983[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_5 (.CI(n16185), .I0(n836_adj_1984[2]), .I1(n206_c), 
            .CO(n16186));
    SB_LUT4 Q_15__I_0_add_564_4_lut (.I0(GND_net), .I1(n836_adj_1984[1]), 
            .I2(n157), .I3(n16184), .O(n835_adj_1983[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_4 (.CI(n16184), .I0(n836_adj_1984[1]), .I1(n157), 
            .CO(n16185));
    SB_LUT4 Q_15__I_0_add_564_3_lut (.I0(GND_net), .I1(n836_adj_1984[0]), 
            .I2(n108), .I3(n16183), .O(n835_adj_1983[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_3 (.CI(n16183), .I0(n836_adj_1984[0]), .I1(n108), 
            .CO(n16184));
    SB_LUT4 Q_15__I_0_add_564_2_lut (.I0(GND_net), .I1(n14), .I2(n59), 
            .I3(GND_net), .O(n835_adj_1983[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_564_2 (.CI(GND_net), .I0(n14), .I1(n59), .CO(n16183));
    SB_LUT4 Q_15__I_0_add_565_16_lut (.I0(GND_net), .I1(n837_adj_1985[13]), 
            .I2(n753), .I3(n16181), .O(n836_adj_1984[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_16 (.CI(n16181), .I0(n837_adj_1985[13]), 
            .I1(n753), .CO(n755_adj_1464));
    SB_LUT4 Q_15__I_0_add_565_15_lut (.I0(GND_net), .I1(n837_adj_1985[12]), 
            .I2(n699), .I3(n16180), .O(n836_adj_1984[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_15 (.CI(n16180), .I0(n837_adj_1985[12]), 
            .I1(n699), .CO(n16181));
    SB_LUT4 Q_15__I_0_add_565_14_lut (.I0(GND_net), .I1(n837_adj_1985[11]), 
            .I2(n650), .I3(n16179), .O(n836_adj_1984[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_14 (.CI(n16179), .I0(n837_adj_1985[11]), 
            .I1(n650), .CO(n16180));
    SB_LUT4 Q_15__I_0_add_565_13_lut (.I0(GND_net), .I1(n837_adj_1985[10]), 
            .I2(n601), .I3(n16178), .O(n836_adj_1984[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_13 (.CI(n16178), .I0(n837_adj_1985[10]), 
            .I1(n601), .CO(n16179));
    SB_LUT4 Q_15__I_0_add_565_12_lut (.I0(GND_net), .I1(n837_adj_1985[9]), 
            .I2(n552), .I3(n16177), .O(n836_adj_1984[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_12 (.CI(n16177), .I0(n837_adj_1985[9]), .I1(n552), 
            .CO(n16178));
    SB_LUT4 Q_15__I_0_add_565_11_lut (.I0(GND_net), .I1(n837_adj_1985[8]), 
            .I2(n503), .I3(n16176), .O(n836_adj_1984[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_11 (.CI(n16176), .I0(n837_adj_1985[8]), .I1(n503), 
            .CO(n16177));
    SB_LUT4 Q_15__I_0_add_565_10_lut (.I0(GND_net), .I1(n837_adj_1985[7]), 
            .I2(n454), .I3(n16175), .O(n836_adj_1984[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_10 (.CI(n16175), .I0(n837_adj_1985[7]), .I1(n454), 
            .CO(n16176));
    SB_LUT4 Q_15__I_0_add_565_9_lut (.I0(GND_net), .I1(n837_adj_1985[6]), 
            .I2(n405_adj_225), .I3(n16174), .O(n836_adj_1984[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_9 (.CI(n16174), .I0(n837_adj_1985[6]), .I1(n405_adj_225), 
            .CO(n16175));
    SB_LUT4 Q_15__I_0_add_565_8_lut (.I0(GND_net), .I1(n837_adj_1985[5]), 
            .I2(n356), .I3(n16173), .O(n836_adj_1984[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_8 (.CI(n16173), .I0(n837_adj_1985[5]), .I1(n356), 
            .CO(n16174));
    SB_LUT4 Q_15__I_0_add_565_7_lut (.I0(GND_net), .I1(n837_adj_1985[4]), 
            .I2(n307), .I3(n16172), .O(n836_adj_1984[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_7 (.CI(n16172), .I0(n837_adj_1985[4]), .I1(n307), 
            .CO(n16173));
    SB_LUT4 Q_15__I_0_add_565_6_lut (.I0(GND_net), .I1(n837_adj_1985[3]), 
            .I2(n258), .I3(n16171), .O(n836_adj_1984[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_6 (.CI(n16171), .I0(n837_adj_1985[3]), .I1(n258), 
            .CO(n16172));
    SB_LUT4 Q_15__I_0_add_565_5_lut (.I0(GND_net), .I1(n837_adj_1985[2]), 
            .I2(n209_c), .I3(n16170), .O(n836_adj_1984[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_5 (.CI(n16170), .I0(n837_adj_1985[2]), .I1(n209_c), 
            .CO(n16171));
    SB_LUT4 Q_15__I_0_add_565_4_lut (.I0(GND_net), .I1(n837_adj_1985[1]), 
            .I2(n160), .I3(n16169), .O(n836_adj_1984[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_4 (.CI(n16169), .I0(n837_adj_1985[1]), .I1(n160), 
            .CO(n16170));
    SB_LUT4 Q_15__I_0_add_565_3_lut (.I0(GND_net), .I1(n837_adj_1985[0]), 
            .I2(n111_adj_226), .I3(n16168), .O(n836_adj_1984[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_3 (.CI(n16168), .I0(n837_adj_1985[0]), .I1(n111_adj_226), 
            .CO(n16169));
    SB_LUT4 Q_15__I_0_add_565_2_lut (.I0(GND_net), .I1(n17), .I2(n62), 
            .I3(GND_net), .O(n836_adj_1984[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_565_2 (.CI(GND_net), .I0(n17), .I1(n62), .CO(n16168));
    SB_LUT4 Q_15__I_0_add_566_16_lut (.I0(GND_net), .I1(n838_adj_1986[13]), 
            .I2(n757), .I3(n16166), .O(n837_adj_1985[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_16 (.CI(n16166), .I0(n838_adj_1986[13]), 
            .I1(n757), .CO(n759_adj_1482));
    SB_LUT4 Q_15__I_0_add_566_15_lut (.I0(GND_net), .I1(n838_adj_1986[12]), 
            .I2(n702), .I3(n16165), .O(n837_adj_1985[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_15 (.CI(n16165), .I0(n838_adj_1986[12]), 
            .I1(n702), .CO(n16166));
    SB_LUT4 Q_15__I_0_add_566_14_lut (.I0(GND_net), .I1(n838_adj_1986[11]), 
            .I2(n653), .I3(n16164), .O(n837_adj_1985[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_14 (.CI(n16164), .I0(n838_adj_1986[11]), 
            .I1(n653), .CO(n16165));
    SB_LUT4 Q_15__I_0_add_566_13_lut (.I0(GND_net), .I1(n838_adj_1986[10]), 
            .I2(n604), .I3(n16163), .O(n837_adj_1985[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_13 (.CI(n16163), .I0(n838_adj_1986[10]), 
            .I1(n604), .CO(n16164));
    SB_LUT4 Q_15__I_0_add_566_12_lut (.I0(GND_net), .I1(n838_adj_1986[9]), 
            .I2(n555), .I3(n16162), .O(n837_adj_1985[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_12 (.CI(n16162), .I0(n838_adj_1986[9]), .I1(n555), 
            .CO(n16163));
    SB_LUT4 Q_15__I_0_add_566_11_lut (.I0(GND_net), .I1(n838_adj_1986[8]), 
            .I2(n506), .I3(n16161), .O(n837_adj_1985[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_11 (.CI(n16161), .I0(n838_adj_1986[8]), .I1(n506), 
            .CO(n16162));
    SB_LUT4 Q_15__I_0_add_566_10_lut (.I0(GND_net), .I1(n838_adj_1986[7]), 
            .I2(n457), .I3(n16160), .O(n837_adj_1985[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_10 (.CI(n16160), .I0(n838_adj_1986[7]), .I1(n457), 
            .CO(n16161));
    SB_LUT4 Q_15__I_0_add_566_9_lut (.I0(GND_net), .I1(n838_adj_1986[6]), 
            .I2(n408), .I3(n16159), .O(n837_adj_1985[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_9 (.CI(n16159), .I0(n838_adj_1986[6]), .I1(n408), 
            .CO(n16160));
    SB_LUT4 Q_15__I_0_add_566_8_lut (.I0(GND_net), .I1(n838_adj_1986[5]), 
            .I2(n359), .I3(n16158), .O(n837_adj_1985[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_8 (.CI(n16158), .I0(n838_adj_1986[5]), .I1(n359), 
            .CO(n16159));
    SB_LUT4 Q_15__I_0_add_566_7_lut (.I0(GND_net), .I1(n838_adj_1986[4]), 
            .I2(n310), .I3(n16157), .O(n837_adj_1985[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_7 (.CI(n16157), .I0(n838_adj_1986[4]), .I1(n310), 
            .CO(n16158));
    SB_LUT4 Q_15__I_0_add_566_6_lut (.I0(GND_net), .I1(n838_adj_1986[3]), 
            .I2(n261), .I3(n16156), .O(n837_adj_1985[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_6 (.CI(n16156), .I0(n838_adj_1986[3]), .I1(n261), 
            .CO(n16157));
    SB_LUT4 Q_15__I_0_add_566_5_lut (.I0(GND_net), .I1(n838_adj_1986[2]), 
            .I2(n212_c), .I3(n16155), .O(n837_adj_1985[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_5 (.CI(n16155), .I0(n838_adj_1986[2]), .I1(n212_c), 
            .CO(n16156));
    SB_LUT4 Q_15__I_0_add_566_4_lut (.I0(GND_net), .I1(n838_adj_1986[1]), 
            .I2(n163), .I3(n16154), .O(n837_adj_1985[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_4 (.CI(n16154), .I0(n838_adj_1986[1]), .I1(n163), 
            .CO(n16155));
    SB_LUT4 Q_15__I_0_add_566_3_lut (.I0(GND_net), .I1(n838_adj_1986[0]), 
            .I2(n114_adj_227), .I3(n16153), .O(n837_adj_1985[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_3 (.CI(n16153), .I0(n838_adj_1986[0]), .I1(n114_adj_227), 
            .CO(n16154));
    SB_LUT4 Q_15__I_0_add_566_2_lut (.I0(GND_net), .I1(n20_adj_228), .I2(n65_adj_229), 
            .I3(GND_net), .O(n837_adj_1985[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_566_2 (.CI(GND_net), .I0(n20_adj_228), .I1(n65_adj_229), 
            .CO(n16153));
    SB_LUT4 Q_15__I_0_add_567_16_lut (.I0(GND_net), .I1(n839_adj_1987[13]), 
            .I2(n761), .I3(n16151), .O(n838_adj_1986[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_16 (.CI(n16151), .I0(n839_adj_1987[13]), 
            .I1(n761), .CO(n763_adj_1502));
    SB_LUT4 Q_15__I_0_add_567_15_lut (.I0(GND_net), .I1(n839_adj_1987[12]), 
            .I2(n705), .I3(n16150), .O(n838_adj_1986[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_15 (.CI(n16150), .I0(n839_adj_1987[12]), 
            .I1(n705), .CO(n16151));
    SB_LUT4 Q_15__I_0_add_567_14_lut (.I0(GND_net), .I1(n839_adj_1987[11]), 
            .I2(n656), .I3(n16149), .O(n838_adj_1986[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_14 (.CI(n16149), .I0(n839_adj_1987[11]), 
            .I1(n656), .CO(n16150));
    SB_LUT4 Q_15__I_0_add_567_13_lut (.I0(GND_net), .I1(n839_adj_1987[10]), 
            .I2(n607), .I3(n16148), .O(n838_adj_1986[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_13 (.CI(n16148), .I0(n839_adj_1987[10]), 
            .I1(n607), .CO(n16149));
    SB_LUT4 Q_15__I_0_add_567_12_lut (.I0(GND_net), .I1(n839_adj_1987[9]), 
            .I2(n558), .I3(n16147), .O(n838_adj_1986[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_12 (.CI(n16147), .I0(n839_adj_1987[9]), .I1(n558), 
            .CO(n16148));
    SB_LUT4 Q_15__I_0_add_567_11_lut (.I0(GND_net), .I1(n839_adj_1987[8]), 
            .I2(n509), .I3(n16146), .O(n838_adj_1986[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_11 (.CI(n16146), .I0(n839_adj_1987[8]), .I1(n509), 
            .CO(n16147));
    SB_LUT4 Q_15__I_0_add_567_10_lut (.I0(GND_net), .I1(n839_adj_1987[7]), 
            .I2(n460), .I3(n16145), .O(n838_adj_1986[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_10 (.CI(n16145), .I0(n839_adj_1987[7]), .I1(n460), 
            .CO(n16146));
    SB_LUT4 Q_15__I_0_add_567_9_lut (.I0(GND_net), .I1(n839_adj_1987[6]), 
            .I2(n411), .I3(n16144), .O(n838_adj_1986[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_9 (.CI(n16144), .I0(n839_adj_1987[6]), .I1(n411), 
            .CO(n16145));
    SB_LUT4 Q_15__I_0_add_567_8_lut (.I0(GND_net), .I1(n839_adj_1987[5]), 
            .I2(n362), .I3(n16143), .O(n838_adj_1986[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_8 (.CI(n16143), .I0(n839_adj_1987[5]), .I1(n362), 
            .CO(n16144));
    SB_LUT4 Q_15__I_0_add_567_7_lut (.I0(GND_net), .I1(n839_adj_1987[4]), 
            .I2(n313_adj_1513), .I3(n16142), .O(n838_adj_1986[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_7 (.CI(n16142), .I0(n839_adj_1987[4]), .I1(n313_adj_1513), 
            .CO(n16143));
    SB_LUT4 Q_15__I_0_add_567_6_lut (.I0(GND_net), .I1(n839_adj_1987[3]), 
            .I2(n264_adj_230), .I3(n16141), .O(n838_adj_1986[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_6 (.CI(n16141), .I0(n839_adj_1987[3]), .I1(n264_adj_230), 
            .CO(n16142));
    SB_LUT4 Q_15__I_0_add_567_5_lut (.I0(GND_net), .I1(n839_adj_1987[2]), 
            .I2(n215_adj_1517), .I3(n16140), .O(n838_adj_1986[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_5 (.CI(n16140), .I0(n839_adj_1987[2]), .I1(n215_adj_1517), 
            .CO(n16141));
    SB_LUT4 Q_15__I_0_add_567_4_lut (.I0(GND_net), .I1(n839_adj_1987[1]), 
            .I2(n166_adj_1519), .I3(n16139), .O(n838_adj_1986[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_4 (.CI(n16139), .I0(n839_adj_1987[1]), .I1(n166_adj_1519), 
            .CO(n16140));
    SB_LUT4 Q_15__I_0_add_567_3_lut (.I0(GND_net), .I1(n839_adj_1987[0]), 
            .I2(n117), .I3(n16138), .O(n838_adj_1986[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_3 (.CI(n16138), .I0(n839_adj_1987[0]), .I1(n117), 
            .CO(n16139));
    SB_LUT4 Q_15__I_0_add_567_2_lut (.I0(GND_net), .I1(n23), .I2(n68), 
            .I3(GND_net), .O(n838_adj_1986[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_567_2 (.CI(GND_net), .I0(n23), .I1(n68), .CO(n16138));
    SB_LUT4 Q_15__I_0_add_568_16_lut (.I0(GND_net), .I1(n840_adj_1988[13]), 
            .I2(n765), .I3(n16136), .O(n839_adj_1987[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_16 (.CI(n16136), .I0(n840_adj_1988[13]), 
            .I1(n765), .CO(n767_adj_1523));
    SB_LUT4 Q_15__I_0_add_568_15_lut (.I0(GND_net), .I1(n840_adj_1988[12]), 
            .I2(n708_adj_1525), .I3(n16135), .O(n839_adj_1987[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_15 (.CI(n16135), .I0(n840_adj_1988[12]), 
            .I1(n708_adj_1525), .CO(n16136));
    SB_LUT4 Q_15__I_0_add_568_14_lut (.I0(GND_net), .I1(n840_adj_1988[11]), 
            .I2(n659_adj_1527), .I3(n16134), .O(n839_adj_1987[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_14 (.CI(n16134), .I0(n840_adj_1988[11]), 
            .I1(n659_adj_1527), .CO(n16135));
    SB_LUT4 Q_15__I_0_add_568_13_lut (.I0(GND_net), .I1(n840_adj_1988[10]), 
            .I2(n610_adj_231), .I3(n16133), .O(n839_adj_1987[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_13 (.CI(n16133), .I0(n840_adj_1988[10]), 
            .I1(n610_adj_231), .CO(n16134));
    SB_LUT4 Q_15__I_0_add_568_12_lut (.I0(GND_net), .I1(n840_adj_1988[9]), 
            .I2(n561), .I3(n16132), .O(n839_adj_1987[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_12 (.CI(n16132), .I0(n840_adj_1988[9]), .I1(n561), 
            .CO(n16133));
    SB_LUT4 Q_15__I_0_add_568_11_lut (.I0(GND_net), .I1(n840_adj_1988[8]), 
            .I2(n512_adj_1533), .I3(n16131), .O(n839_adj_1987[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_11 (.CI(n16131), .I0(n840_adj_1988[8]), .I1(n512_adj_1533), 
            .CO(n16132));
    SB_LUT4 Q_15__I_0_add_568_10_lut (.I0(GND_net), .I1(n840_adj_1988[7]), 
            .I2(n463_adj_1535), .I3(n16130), .O(n839_adj_1987[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_10 (.CI(n16130), .I0(n840_adj_1988[7]), .I1(n463_adj_1535), 
            .CO(n16131));
    SB_LUT4 Q_15__I_0_add_568_9_lut (.I0(GND_net), .I1(n840_adj_1988[6]), 
            .I2(n414_adj_232), .I3(n16129), .O(n839_adj_1987[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_9 (.CI(n16129), .I0(n840_adj_1988[6]), .I1(n414_adj_232), 
            .CO(n16130));
    SB_LUT4 Q_15__I_0_add_568_8_lut (.I0(GND_net), .I1(n840_adj_1988[5]), 
            .I2(n365_adj_1539), .I3(n16128), .O(n839_adj_1987[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_8 (.CI(n16128), .I0(n840_adj_1988[5]), .I1(n365_adj_1539), 
            .CO(n16129));
    SB_LUT4 Q_15__I_0_add_568_7_lut (.I0(GND_net), .I1(n840_adj_1988[4]), 
            .I2(n316_adj_1541), .I3(n16127), .O(n839_adj_1987[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_11_lut (.I0(GND_net), .I1(n839_adj_1951[8]), 
            .I2(n509_adj_1542), .I3(n16803), .O(n838[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_7 (.CI(n16127), .I0(n840_adj_1988[4]), .I1(n316_adj_1541), 
            .CO(n16128));
    SB_LUT4 Q_15__I_0_add_568_6_lut (.I0(GND_net), .I1(n840_adj_1988[3]), 
            .I2(n267_adj_233), .I3(n16126), .O(n839_adj_1987[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_6 (.CI(n16126), .I0(n840_adj_1988[3]), .I1(n267_adj_233), 
            .CO(n16127));
    SB_CARRY D_15__I_0_10_add_567_11 (.CI(n16803), .I0(n839_adj_1951[8]), 
            .I1(n509_adj_1542), .CO(n16804));
    SB_LUT4 Q_15__I_0_add_568_5_lut (.I0(GND_net), .I1(n840_adj_1988[2]), 
            .I2(n218_adj_1546), .I3(n16125), .O(n839_adj_1987[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_16_lut (.I0(GND_net), .I1(n839_adj_1951[13]), 
            .I2(n761_adj_234), .I3(n16808), .O(n838[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_5 (.CI(n16125), .I0(n840_adj_1988[2]), .I1(n218_adj_1546), 
            .CO(n16126));
    SB_LUT4 Q_15__I_0_add_568_4_lut (.I0(GND_net), .I1(n840_adj_1988[1]), 
            .I2(n169_adj_1550), .I3(n16124), .O(n839_adj_1987[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_4 (.CI(n16124), .I0(n840_adj_1988[1]), .I1(n169_adj_1550), 
            .CO(n16125));
    SB_LUT4 Q_15__I_0_add_568_3_lut (.I0(GND_net), .I1(n840_adj_1988[0]), 
            .I2(n120_adj_235), .I3(n16123), .O(n839_adj_1987[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_3 (.CI(n16123), .I0(n840_adj_1988[0]), .I1(n120_adj_235), 
            .CO(n16124));
    SB_LUT4 Q_15__I_0_add_568_2_lut (.I0(GND_net), .I1(n26_adj_236), .I2(n71_adj_237), 
            .I3(GND_net), .O(n839_adj_1987[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_566_10_lut (.I0(GND_net), .I1(n838[7]), .I2(n457_adj_1557), 
            .I3(n16817), .O(n837[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_568_2 (.CI(GND_net), .I0(n26_adj_236), .I1(n71_adj_237), 
            .CO(n16123));
    SB_LUT4 Q_15__I_0_add_569_16_lut (.I0(GND_net), .I1(n841_adj_1989[13]), 
            .I2(n769_adj_238), .I3(n16121), .O(n840_adj_1988[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_16 (.CI(n16121), .I0(n841_adj_1989[13]), 
            .I1(n769_adj_238), .CO(n771_adj_1561));
    SB_LUT4 Q_15__I_0_add_569_15_lut (.I0(GND_net), .I1(n841_adj_1989[12]), 
            .I2(n711_adj_1563), .I3(n16120), .O(n840_adj_1988[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_15 (.CI(n16120), .I0(n841_adj_1989[12]), 
            .I1(n711_adj_1563), .CO(n16121));
    SB_LUT4 Q_15__I_0_add_569_14_lut (.I0(GND_net), .I1(n841_adj_1989[11]), 
            .I2(n662_adj_1565), .I3(n16119), .O(n840_adj_1988[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_14 (.CI(n16119), .I0(n841_adj_1989[11]), 
            .I1(n662_adj_1565), .CO(n16120));
    SB_LUT4 Q_15__I_0_add_569_13_lut (.I0(GND_net), .I1(n841_adj_1989[10]), 
            .I2(n613_adj_239), .I3(n16118), .O(n840_adj_1988[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_13 (.CI(n16118), .I0(n841_adj_1989[10]), 
            .I1(n613_adj_239), .CO(n16119));
    SB_LUT4 Q_15__I_0_add_569_12_lut (.I0(GND_net), .I1(n841_adj_1989[9]), 
            .I2(n564), .I3(n16117), .O(n840_adj_1988[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_12 (.CI(n16117), .I0(n841_adj_1989[9]), .I1(n564), 
            .CO(n16118));
    SB_LUT4 Q_15__I_0_add_569_11_lut (.I0(GND_net), .I1(n841_adj_1989[8]), 
            .I2(n515_adj_1571), .I3(n16116), .O(n840_adj_1988[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_11 (.CI(n16116), .I0(n841_adj_1989[8]), .I1(n515_adj_1571), 
            .CO(n16117));
    SB_LUT4 Q_15__I_0_add_569_10_lut (.I0(GND_net), .I1(n841_adj_1989[7]), 
            .I2(n466_adj_1573), .I3(n16115), .O(n840_adj_1988[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_10 (.CI(n16115), .I0(n841_adj_1989[7]), .I1(n466_adj_1573), 
            .CO(n16116));
    SB_LUT4 Q_15__I_0_add_569_9_lut (.I0(GND_net), .I1(n841_adj_1989[6]), 
            .I2(n417_adj_240), .I3(n16114), .O(n840_adj_1988[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_9 (.CI(n16114), .I0(n841_adj_1989[6]), .I1(n417_adj_240), 
            .CO(n16115));
    SB_LUT4 Q_15__I_0_add_569_8_lut (.I0(GND_net), .I1(n841_adj_1989[5]), 
            .I2(n368_adj_1577), .I3(n16113), .O(n840_adj_1988[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_8 (.CI(n16113), .I0(n841_adj_1989[5]), .I1(n368_adj_1577), 
            .CO(n16114));
    SB_CARRY Q_15__I_0_11_add_570_13 (.CI(n16566), .I0(n842[10]), .I1(n625_c), 
            .CO(n16567));
    SB_CARRY D_15__I_0_10_add_575_7 (.CI(n16680), .I0(n293_adj_1386), .I1(n337), 
            .CO(n16681));
    SB_CARRY D_15__I_0_10_add_565_3 (.CI(n16825), .I0(n837[0]), .I1(n111), 
            .CO(n16826));
    SB_LUT4 D_15__I_0_10_add_565_2_lut (.I0(GND_net), .I1(n17_adj_241), 
            .I2(n62_adj_242), .I3(GND_net), .O(n836_adj_1960[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_9 (.CI(n16831), .I0(n837[6]), .I1(n405), 
            .CO(n16832));
    SB_LUT4 D_15__I_0_10_add_565_13_lut (.I0(GND_net), .I1(n837[10]), .I2(n601_adj_243), 
            .I3(n16835), .O(n836_adj_1960[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_570_12_lut (.I0(GND_net), .I1(n842[9]), .I2(n576), 
            .I3(n16565), .O(n841_adj_1952[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_6_lut (.I0(GND_net), .I1(n244_adj_244), 
            .I2(n288), .I3(n16679), .O(n846[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_12 (.CI(n16565), .I0(n842[9]), .I1(n576), 
            .CO(n16566));
    SB_CARRY D_15__I_0_10_add_575_6 (.CI(n16679), .I0(n244_adj_244), .I1(n288), 
            .CO(n16680));
    SB_LUT4 Q_15__I_0_11_add_570_11_lut (.I0(GND_net), .I1(n842[8]), .I2(n527), 
            .I3(n16564), .O(n841_adj_1952[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_5_lut (.I0(GND_net), .I1(n195), .I2(n239), 
            .I3(n16678), .O(n846[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_11 (.CI(n16564), .I0(n842[8]), .I1(n527), 
            .CO(n16565));
    SB_LUT4 sub_66_add_2_30_lut (.I0(GND_net), .I1(Product1_mul_temp[29]), 
            .I2(n1[29]), .I3(n17331), .O(alphaVoltage[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_66_add_2_29_lut (.I0(GND_net), .I1(Product1_mul_temp[29]), 
            .I2(n1[29]), .I3(n17330), .O(alphaVoltage[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_29 (.CI(n17330), .I0(Product1_mul_temp[29]), .I1(n1[29]), 
            .CO(n17331));
    SB_LUT4 sub_66_add_2_28_lut (.I0(GND_net), .I1(Product1_mul_temp[28]), 
            .I2(n1[28]), .I3(n17329), .O(alphaVoltage[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_28 (.CI(n17329), .I0(Product1_mul_temp[28]), .I1(n1[28]), 
            .CO(n17330));
    SB_CARRY D_15__I_0_10_add_564_11 (.CI(n16848), .I0(n836_adj_1960[8]), 
            .I1(n500_adj_1590), .CO(n16849));
    SB_LUT4 D_15__I_0_10_add_564_4_lut (.I0(GND_net), .I1(n836_adj_1960[1]), 
            .I2(n157_adj_1592), .I3(n16841), .O(n835_adj_1961[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_4 (.CI(n16841), .I0(n836_adj_1960[1]), 
            .I1(n157_adj_1592), .CO(n16842));
    SB_LUT4 sub_66_add_2_27_lut (.I0(GND_net), .I1(Product1_mul_temp[27]), 
            .I2(n1[27]), .I3(n17328), .O(alphaVoltage[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_5 (.CI(n16678), .I0(n195), .I1(n239), 
            .CO(n16679));
    SB_CARRY sub_66_add_2_27 (.CI(n17328), .I0(Product1_mul_temp[27]), .I1(n1[27]), 
            .CO(n17329));
    SB_LUT4 sub_66_add_2_26_lut (.I0(GND_net), .I1(Product1_mul_temp[26]), 
            .I2(n1[26]), .I3(n17327), .O(alphaVoltage[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_26 (.CI(n17327), .I0(Product1_mul_temp[26]), .I1(n1[26]), 
            .CO(n17328));
    SB_LUT4 sub_66_add_2_25_lut (.I0(GND_net), .I1(Product1_mul_temp[25]), 
            .I2(n1[25]), .I3(n17326), .O(alphaVoltage[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_25 (.CI(n17326), .I0(Product1_mul_temp[25]), .I1(n1[25]), 
            .CO(n17327));
    SB_CARRY D_15__I_0_10_add_564_10 (.CI(n16847), .I0(n836_adj_1960[7]), 
            .I1(n451_adj_1397), .CO(n16848));
    SB_LUT4 Q_15__I_0_add_569_7_lut (.I0(GND_net), .I1(n841_adj_1989[4]), 
            .I2(n319_adj_1594), .I3(n16112), .O(n840_adj_1988[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_66_add_2_24_lut (.I0(GND_net), .I1(Product1_mul_temp[24]), 
            .I2(n1[24]), .I3(n17325), .O(alphaVoltage[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_7 (.CI(n16112), .I0(n841_adj_1989[4]), .I1(n319_adj_1594), 
            .CO(n16113));
    SB_CARRY D_15__I_0_10_add_566_10 (.CI(n16817), .I0(n838[7]), .I1(n457_adj_1557), 
            .CO(n16818));
    SB_CARRY D_15__I_0_10_add_568_14 (.CI(n16791), .I0(n840_adj_1950[11]), 
            .I1(n659), .CO(n16792));
    SB_LUT4 D_15__I_0_10_add_568_13_lut (.I0(GND_net), .I1(n840_adj_1950[10]), 
            .I2(n610), .I3(n16790), .O(n839_adj_1951[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_24 (.CI(n17325), .I0(Product1_mul_temp[24]), .I1(n1[24]), 
            .CO(n17326));
    SB_LUT4 sub_66_add_2_23_lut (.I0(GND_net), .I1(Product1_mul_temp[23]), 
            .I2(n1[23]), .I3(n17324), .O(alphaVoltage[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_23 (.CI(n17324), .I0(Product1_mul_temp[23]), .I1(n1[23]), 
            .CO(n17325));
    SB_CARRY D_15__I_0_10_add_567_4 (.CI(n16796), .I0(n839_adj_1951[1]), 
            .I1(n166), .CO(n16797));
    SB_LUT4 Q_15__I_0_11_add_570_10_lut (.I0(GND_net), .I1(n842[7]), .I2(n478), 
            .I3(n16563), .O(n841_adj_1952[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_10_lut (.I0(GND_net), .I1(n839_adj_1951[7]), 
            .I2(n460_adj_1598), .I3(n16802), .O(n838[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_16 (.CI(n16808), .I0(n839_adj_1951[13]), 
            .I1(n761_adj_234), .CO(n763));
    SB_LUT4 D_15__I_0_10_add_567_15_lut (.I0(GND_net), .I1(n839_adj_1951[12]), 
            .I2(n705_adj_1600), .I3(n16807), .O(n838[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_66_add_2_22_lut (.I0(GND_net), .I1(Product1_mul_temp[22]), 
            .I2(n1[22]), .I3(n17323), .O(alphaVoltage[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_566_9_lut (.I0(GND_net), .I1(n838[6]), .I2(n408_adj_245), 
            .I3(n16816), .O(n837[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_2 (.CI(GND_net), .I0(n17_adj_241), .I1(n62_adj_242), 
            .CO(n16825));
    SB_LUT4 D_15__I_0_10_add_565_8_lut (.I0(GND_net), .I1(n837[5]), .I2(n356_adj_1605), 
            .I3(n16830), .O(n836_adj_1960[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_8 (.CI(n16830), .I0(n837[5]), .I1(n356_adj_1605), 
            .CO(n16831));
    SB_CARRY sub_66_add_2_22 (.CI(n17323), .I0(Product1_mul_temp[22]), .I1(n1[22]), 
            .CO(n17324));
    SB_CARRY D_15__I_0_10_add_565_13 (.CI(n16835), .I0(n837[10]), .I1(n601_adj_243), 
            .CO(n16836));
    SB_CARRY D_15__I_0_10_add_567_15 (.CI(n16807), .I0(n839_adj_1951[12]), 
            .I1(n705_adj_1600), .CO(n16808));
    SB_LUT4 D_15__I_0_10_add_564_3_lut (.I0(GND_net), .I1(n836_adj_1960[0]), 
            .I2(n108_adj_246), .I3(n16840), .O(n835_adj_1961[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_4_lut (.I0(GND_net), .I1(n146_adj_1608), 
            .I2(n190), .I3(n16677), .O(n846[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_564_9_lut (.I0(GND_net), .I1(n836_adj_1960[6]), 
            .I2(n402_adj_247), .I3(n16846), .O(n835_adj_1961[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_9 (.CI(n16846), .I0(n836_adj_1960[6]), 
            .I1(n402_adj_247), .CO(n16847));
    SB_LUT4 sub_66_add_2_21_lut (.I0(GND_net), .I1(Product1_mul_temp[21]), 
            .I2(n1[21]), .I3(n17322), .O(alphaVoltage[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_9 (.CI(n16816), .I0(n838[6]), .I1(n408_adj_245), 
            .CO(n16817));
    SB_LUT4 Q_15__I_0_add_569_6_lut (.I0(GND_net), .I1(n841_adj_1989[3]), 
            .I2(n270_adj_248), .I3(n16111), .O(n840_adj_1988[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_21 (.CI(n17322), .I0(Product1_mul_temp[21]), .I1(n1[21]), 
            .CO(n17323));
    SB_LUT4 sub_66_add_2_20_lut (.I0(GND_net), .I1(Product1_mul_temp[20]), 
            .I2(n1[20]), .I3(n17321), .O(alphaVoltage[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_6 (.CI(n16111), .I0(n841_adj_1989[3]), .I1(n270_adj_248), 
            .CO(n16112));
    SB_CARRY sub_66_add_2_20 (.CI(n17321), .I0(Product1_mul_temp[20]), .I1(n1[20]), 
            .CO(n17322));
    SB_LUT4 D_15__I_0_10_add_564_14_lut (.I0(GND_net), .I1(n836_adj_1960[11]), 
            .I2(n647_adj_1614), .I3(n16851), .O(n835_adj_1961[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_66_add_2_19_lut (.I0(GND_net), .I1(Product1_mul_temp[19]), 
            .I2(n1[19]), .I3(n17320), .O(alphaVoltage[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_563_9 (.CI(n16861), .I0(n835_adj_1961[6]), 
            .I1(n399), .CO(n16862));
    SB_CARRY sub_66_add_2_19 (.CI(n17320), .I0(Product1_mul_temp[19]), .I1(n1[19]), 
            .CO(n17321));
    SB_CARRY D_15__I_0_10_add_562_2 (.CI(GND_net), .I0(n8), .I1(n53), 
            .CO(n16870));
    SB_CARRY Q_15__I_0_11_add_570_10 (.CI(n16563), .I0(n842[7]), .I1(n478), 
            .CO(n16564));
    SB_LUT4 D_15__I_0_10_add_563_16_lut (.I0(GND_net), .I1(n835_adj_1961[13]), 
            .I2(n745_adj_249), .I3(n16868), .O(n834[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_66_add_2_18_lut (.I0(GND_net), .I1(Product1_mul_temp[18]), 
            .I2(n1[18]), .I3(n17319), .O(alphaVoltage[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_562_11_lut (.I0(GND_net), .I1(n834[8]), .I2(n494_adj_1618), 
            .I3(n16878), .O(n833[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_14 (.CI(n16851), .I0(n836_adj_1960[11]), 
            .I1(n647_adj_1614), .CO(n16852));
    SB_CARRY sub_66_add_2_18 (.CI(n17319), .I0(Product1_mul_temp[18]), .I1(n1[18]), 
            .CO(n17320));
    SB_LUT4 sub_66_add_2_17_lut (.I0(GND_net), .I1(Product1_mul_temp[17]), 
            .I2(n1[17]), .I3(n17318), .O(alphaVoltage[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_17 (.CI(n17318), .I0(Product1_mul_temp[17]), .I1(n1[17]), 
            .CO(n17319));
    SB_CARRY D_15__I_0_10_add_561_7 (.CI(n16889), .I0(n833[4]), .I1(n295_adj_1333), 
            .CO(n16890));
    SB_LUT4 D_15__I_0_10_add_561_15_lut (.I0(GND_net), .I1(n833[12]), .I2(n687_adj_1620), 
            .I3(n16897), .O(Product1_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_15 (.CI(n16897), .I0(n833[12]), .I1(n687_adj_1620), 
            .CO(n16898));
    SB_LUT4 sub_66_add_2_16_lut (.I0(GND_net), .I1(Product1_mul_temp[16]), 
            .I2(n1[16]), .I3(n17317), .O(alphaVoltage[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_564_11_lut (.I0(GND_net), .I1(n836_adj_1960[8]), 
            .I2(n500_adj_1590), .I3(n16848), .O(n835_adj_1961[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_4 (.CI(n16677), .I0(n146_adj_1608), .I1(n190), 
            .CO(n16678));
    SB_CARRY sub_66_add_2_16 (.CI(n17317), .I0(Product1_mul_temp[16]), .I1(n1[16]), 
            .CO(n17318));
    SB_LUT4 sub_66_add_2_15_lut (.I0(GND_net), .I1(Product1_mul_temp[15]), 
            .I2(n1[15]), .I3(n17316), .O(alphaVoltage[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_66_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_8_lut (.I0(GND_net), .I1(n835_adj_1961[5]), 
            .I2(n350_adj_1625), .I3(n16860), .O(n834[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_15 (.CI(n17316), .I0(Product1_mul_temp[15]), .I1(n1[15]), 
            .CO(n17317));
    SB_CARRY sub_66_add_2_14 (.CI(n17315), .I0(Product1_mul_temp[14]), .I1(n1[14]), 
            .CO(n17316));
    SB_LUT4 Q_15__I_0_11_add_570_9_lut (.I0(GND_net), .I1(n842[6]), .I2(n429_c), 
            .I3(n16562), .O(n841_adj_1952[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_13 (.CI(n17314), .I0(Product1_mul_temp[13]), .I1(n1[13]), 
            .CO(n17315));
    SB_CARRY D_15__I_0_10_add_563_8 (.CI(n16860), .I0(n835_adj_1961[5]), 
            .I1(n350_adj_1625), .CO(n16861));
    SB_LUT4 D_15__I_0_10_add_563_7_lut (.I0(GND_net), .I1(n835_adj_1961[4]), 
            .I2(n301_adj_1629), .I3(n16859), .O(n834[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_12 (.CI(n17313), .I0(Product1_mul_temp[12]), .I1(n1[12]), 
            .CO(n17314));
    SB_CARRY sub_66_add_2_11 (.CI(n17312), .I0(Product1_mul_temp[11]), .I1(n1[11]), 
            .CO(n17313));
    SB_CARRY sub_66_add_2_10 (.CI(n17311), .I0(Product1_mul_temp[10]), .I1(n1[10]), 
            .CO(n17312));
    SB_CARRY sub_66_add_2_9 (.CI(n17310), .I0(Product1_mul_temp[9]), .I1(n1[9]), 
            .CO(n17311));
    SB_CARRY sub_66_add_2_8 (.CI(n17309), .I0(Product1_mul_temp[8]), .I1(n1[8]), 
            .CO(n17310));
    SB_CARRY sub_66_add_2_7 (.CI(n17308), .I0(Product1_mul_temp[7]), .I1(n1[7]), 
            .CO(n17309));
    SB_CARRY sub_66_add_2_6 (.CI(n17307), .I0(Product1_mul_temp[6]), .I1(n1[6]), 
            .CO(n17308));
    SB_CARRY D_15__I_0_10_add_563_7 (.CI(n16859), .I0(n835_adj_1961[4]), 
            .I1(n301_adj_1629), .CO(n16860));
    SB_CARRY D_15__I_0_10_add_563_16 (.CI(n16868), .I0(n835_adj_1961[13]), 
            .I1(n745_adj_249), .CO(n747));
    SB_CARRY sub_66_add_2_5 (.CI(n17306), .I0(Product1_mul_temp[5]), .I1(n1[5]), 
            .CO(n17307));
    SB_CARRY D_15__I_0_10_add_562_11 (.CI(n16878), .I0(n834[8]), .I1(n494_adj_1618), 
            .CO(n16879));
    SB_CARRY sub_66_add_2_4 (.CI(n17305), .I0(Product1_mul_temp[4]), .I1(n1[4]), 
            .CO(n17306));
    SB_LUT4 D_15__I_0_10_add_575_3_lut (.I0(GND_net), .I1(n97_adj_1633), 
            .I2(n141), .I3(n16676), .O(n846[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_6_lut (.I0(GND_net), .I1(n833[3]), .I2(n246_adj_250), 
            .I3(n16888), .O(Product1_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_66_add_2_3 (.CI(n17304), .I0(Product1_mul_temp[3]), .I1(n1[3]), 
            .CO(n17305));
    SB_CARRY sub_66_add_2_2 (.CI(VCC_net), .I0(Product1_mul_temp[2]), .I1(n1[2]), 
            .CO(n17304));
    SB_LUT4 Q_15__I_0_add_569_5_lut (.I0(GND_net), .I1(n841_adj_1989[2]), 
            .I2(n221_adj_1638), .I3(n16110), .O(n840_adj_1988[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_5 (.CI(n16110), .I0(n841_adj_1989[2]), .I1(n221_adj_1638), 
            .CO(n16111));
    SB_CARRY Q_15__I_0_11_add_570_9 (.CI(n16562), .I0(n842[6]), .I1(n429_c), 
            .CO(n16563));
    SB_LUT4 Q_15__I_0_add_569_4_lut (.I0(GND_net), .I1(n841_adj_1989[1]), 
            .I2(n172_adj_1640), .I3(n16109), .O(n840_adj_1988[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_4 (.CI(n16109), .I0(n841_adj_1989[1]), .I1(n172_adj_1640), 
            .CO(n16110));
    SB_LUT4 Q_15__I_0_add_569_3_lut (.I0(GND_net), .I1(n841_adj_1989[0]), 
            .I2(n123_adj_251), .I3(n16108), .O(n840_adj_1988[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_3_lut (.I0(GND_net), .I1(n839_adj_1951[0]), 
            .I2(n117_adj_252), .I3(n16795), .O(n838[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_3 (.CI(n16795), .I0(n839_adj_1951[0]), 
            .I1(n117_adj_252), .CO(n16796));
    SB_CARRY D_15__I_0_10_add_567_10 (.CI(n16802), .I0(n839_adj_1951[7]), 
            .I1(n460_adj_1598), .CO(n16803));
    SB_CARRY D_15__I_0_10_add_561_6 (.CI(n16888), .I0(n833[3]), .I1(n246_adj_250), 
            .CO(n16889));
    SB_LUT4 D_15__I_0_10_add_567_14_lut (.I0(GND_net), .I1(n839_adj_1951[11]), 
            .I2(n656_adj_1646), .I3(n16806), .O(n838[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_3 (.CI(n16676), .I0(n97_adj_1633), .I1(n141), 
            .CO(n16677));
    SB_LUT4 D_15__I_0_10_add_566_8_lut (.I0(GND_net), .I1(n838[5]), .I2(n359_adj_1648), 
            .I3(n16815), .O(n837[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_14_lut (.I0(GND_net), .I1(n833[11]), .I2(n638_adj_1649), 
            .I3(n16896), .O(Product1_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_8 (.CI(n16815), .I0(n838[5]), .I1(n359_adj_1648), 
            .CO(n16816));
    SB_LUT4 D_15__I_0_10_add_566_16_lut (.I0(GND_net), .I1(n838[13]), .I2(n757_adj_253), 
            .I3(n16823), .O(n837[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_565_7_lut (.I0(GND_net), .I1(n837[4]), .I2(n307_adj_1653), 
            .I3(n16829), .O(n836_adj_1960[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_565_12_lut (.I0(GND_net), .I1(n837[9]), .I2(n552_adj_1654), 
            .I3(n16834), .O(n836_adj_1960[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_12 (.CI(n16834), .I0(n837[9]), .I1(n552_adj_1654), 
            .CO(n16835));
    SB_CARRY D_15__I_0_10_add_564_3 (.CI(n16840), .I0(n836_adj_1960[0]), 
            .I1(n108_adj_246), .CO(n16841));
    SB_LUT4 D_15__I_0_10_add_564_8_lut (.I0(GND_net), .I1(n836_adj_1960[5]), 
            .I2(n353_adj_1655), .I3(n16845), .O(n835_adj_1961[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_15_lut (.I0(GND_net), .I1(n835_adj_1961[12]), 
            .I2(n693_adj_1657), .I3(n16867), .O(n834[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_2_lut (.I0(GND_net), .I1(n23_adj_254), 
            .I2(n68_adj_255), .I3(GND_net), .O(n838[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_570_8_lut (.I0(GND_net), .I1(n842[5]), .I2(n380), 
            .I3(n16561), .O(n841_adj_1952[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_566_7_lut (.I0(GND_net), .I1(n838[4]), .I2(n310_adj_1660), 
            .I3(n16814), .O(n837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_3 (.CI(n16108), .I0(n841_adj_1989[0]), .I1(n123_adj_251), 
            .CO(n16109));
    SB_CARRY D_15__I_0_10_add_564_12 (.CI(n16849), .I0(n836_adj_1960[9]), 
            .I1(n549_adj_1662), .CO(n16850));
    SB_LUT4 D_15__I_0_10_add_572_10_lut (.I0(GND_net), .I1(n844_adj_1959[7]), 
            .I2(n475), .I3(n16727), .O(n843_adj_1956[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_6_lut (.I0(GND_net), .I1(n835_adj_1961[3]), 
            .I2(n252_adj_256), .I3(n16858), .O(n834[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_563_15 (.CI(n16867), .I0(n835_adj_1961[12]), 
            .I1(n693_adj_1657), .CO(n16868));
    SB_LUT4 D_15__I_0_10_add_562_10_lut (.I0(GND_net), .I1(n834[7]), .I2(n445_adj_1667), 
            .I3(n16877), .O(n833[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_10 (.CI(n16877), .I0(n834[7]), .I1(n445_adj_1667), 
            .CO(n16878));
    SB_LUT4 D_15__I_0_10_add_562_9_lut (.I0(GND_net), .I1(n834[6]), .I2(n396_adj_257), 
            .I3(n16876), .O(n833[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_575_2_lut (.I0(GND_net), .I1(n48_adj_1670), 
            .I2(n92), .I3(GND_net), .O(n846[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_575_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_5_lut (.I0(GND_net), .I1(n833[2]), .I2(n197), 
            .I3(n16887), .O(Product1_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_14 (.CI(n16896), .I0(n833[11]), .I1(n638_adj_1649), 
            .CO(n16897));
    SB_CARRY D_15__I_0_10_add_561_5 (.CI(n16887), .I0(n833[2]), .I1(n197), 
            .CO(n16888));
    SB_CARRY Q_15__I_0_11_add_570_8 (.CI(n16561), .I0(n842[5]), .I1(n380), 
            .CO(n16562));
    SB_LUT4 D_15__I_0_10_add_561_4_lut (.I0(GND_net), .I1(n833[1]), .I2(n148_adj_1673), 
            .I3(n16886), .O(Product1_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_575_2 (.CI(GND_net), .I0(n48_adj_1670), .I1(n92), 
            .CO(n16676));
    SB_LUT4 Q_15__I_0_11_add_570_7_lut (.I0(GND_net), .I1(n842[4]), .I2(n331), 
            .I3(n16560), .O(n841_adj_1952[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_16_lut (.I0(GND_net), .I1(n835[13]), .I2(n793), 
            .I3(n16674), .O(n834_adj_1976[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_add_569_2_lut (.I0(GND_net), .I1(n29_adj_258), .I2(n74_adj_259), 
            .I3(GND_net), .O(n840_adj_1988[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_569_2 (.CI(GND_net), .I0(n29_adj_258), .I1(n74_adj_259), 
            .CO(n16108));
    SB_LUT4 Q_15__I_0_add_570_16_lut (.I0(GND_net), .I1(n842_adj_1990[13]), 
            .I2(n773_adj_260), .I3(n16106), .O(n841_adj_1989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_16 (.CI(n16106), .I0(n842_adj_1990[13]), 
            .I1(n773_adj_260), .CO(n775_adj_1680));
    SB_LUT4 i7334_2_lut (.I0(n833_adj_1964[13]), .I1(\dVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n832_adj_1979[14]));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam i7334_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Q_15__I_0_add_570_15_lut (.I0(GND_net), .I1(n842_adj_1990[12]), 
            .I2(n714_adj_1682), .I3(n16105), .O(n841_adj_1989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_15 (.CI(n16105), .I0(n842_adj_1990[12]), 
            .I1(n714_adj_1682), .CO(n16106));
    SB_LUT4 D_15__I_0_10_i228_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n337));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_add_570_14_lut (.I0(GND_net), .I1(n842_adj_1990[11]), 
            .I2(n665_adj_1684), .I3(n16104), .O(n841_adj_1989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_14 (.CI(n16104), .I0(n842_adj_1990[11]), 
            .I1(n665_adj_1684), .CO(n16105));
    SB_LUT4 Q_15__I_0_add_570_13_lut (.I0(GND_net), .I1(n842_adj_1990[10]), 
            .I2(n616_adj_261), .I3(n16103), .O(n841_adj_1989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_13 (.CI(n16103), .I0(n842_adj_1990[10]), 
            .I1(n616_adj_261), .CO(n16104));
    SB_LUT4 Q_15__I_0_add_570_12_lut (.I0(GND_net), .I1(n842_adj_1990[9]), 
            .I2(n567), .I3(n16102), .O(n841_adj_1989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_12 (.CI(n16102), .I0(n842_adj_1990[9]), .I1(n567), 
            .CO(n16103));
    SB_LUT4 D_15__I_0_10_i198_2_lut (.I0(\dVoltage[5] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_1386));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i198_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_add_570_11_lut (.I0(GND_net), .I1(n842_adj_1990[8]), 
            .I2(n518_adj_1690), .I3(n16101), .O(n841_adj_1989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_11 (.CI(n16101), .I0(n842_adj_1990[8]), .I1(n518_adj_1690), 
            .CO(n16102));
    SB_LUT4 Q_15__I_0_add_570_10_lut (.I0(GND_net), .I1(n842_adj_1990[7]), 
            .I2(n469_adj_1692), .I3(n16100), .O(n841_adj_1989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_10 (.CI(n16100), .I0(n842_adj_1990[7]), .I1(n469_adj_1692), 
            .CO(n16101));
    SB_LUT4 Q_15__I_0_add_570_9_lut (.I0(GND_net), .I1(n842_adj_1990[6]), 
            .I2(n420_adj_262), .I3(n16099), .O(n841_adj_1989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_9 (.CI(n16099), .I0(n842_adj_1990[6]), .I1(n420_adj_262), 
            .CO(n16100));
    SB_LUT4 Q_15__I_0_add_570_8_lut (.I0(GND_net), .I1(n842_adj_1990[5]), 
            .I2(n371_adj_1696), .I3(n16098), .O(n841_adj_1989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_8 (.CI(n16098), .I0(n842_adj_1990[5]), .I1(n371_adj_1696), 
            .CO(n16099));
    SB_LUT4 Q_15__I_0_add_570_7_lut (.I0(GND_net), .I1(n842_adj_1990[4]), 
            .I2(n322_adj_1698), .I3(n16097), .O(n841_adj_1989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_7 (.CI(n16097), .I0(n842_adj_1990[4]), .I1(n322_adj_1698), 
            .CO(n16098));
    SB_LUT4 Q_15__I_0_add_570_6_lut (.I0(GND_net), .I1(n842_adj_1990[3]), 
            .I2(n273_adj_263), .I3(n16096), .O(n841_adj_1989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_6 (.CI(n16096), .I0(n842_adj_1990[3]), .I1(n273_adj_263), 
            .CO(n16097));
    SB_LUT4 Q_15__I_0_add_570_5_lut (.I0(GND_net), .I1(n842_adj_1990[2]), 
            .I2(n224_adj_1702), .I3(n16095), .O(n841_adj_1989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_5 (.CI(n16095), .I0(n842_adj_1990[2]), .I1(n224_adj_1702), 
            .CO(n16096));
    SB_LUT4 Q_15__I_0_add_570_4_lut (.I0(GND_net), .I1(n842_adj_1990[1]), 
            .I2(n175_adj_1704), .I3(n16094), .O(n841_adj_1989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_4 (.CI(n16094), .I0(n842_adj_1990[1]), .I1(n175_adj_1704), 
            .CO(n16095));
    SB_LUT4 Q_15__I_0_11_i468_2_lut (.I0(\qVoltage[14] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n723));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_add_570_3_lut (.I0(GND_net), .I1(n842_adj_1990[0]), 
            .I2(n126_adj_264), .I3(n16093), .O(n841_adj_1989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_3 (.CI(n16093), .I0(n842_adj_1990[0]), .I1(n126_adj_264), 
            .CO(n16094));
    SB_LUT4 Q_15__I_0_add_570_2_lut (.I0(GND_net), .I1(n32_adj_265), .I2(n77_adj_266), 
            .I3(GND_net), .O(n841_adj_1989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_570_2 (.CI(GND_net), .I0(n32_adj_265), .I1(n77_adj_266), 
            .CO(n16093));
    SB_LUT4 Q_15__I_0_add_571_16_lut (.I0(GND_net), .I1(n843_adj_1991[13]), 
            .I2(n777_adj_267), .I3(n16091), .O(n842_adj_1990[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_16 (.CI(n16091), .I0(n843_adj_1991[13]), 
            .I1(n777_adj_267), .CO(n779_adj_1712));
    SB_LUT4 Q_15__I_0_add_571_15_lut (.I0(GND_net), .I1(n843_adj_1991[12]), 
            .I2(n717_adj_1714), .I3(n16090), .O(n842_adj_1990[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_15 (.CI(n16090), .I0(n843_adj_1991[12]), 
            .I1(n717_adj_1714), .CO(n16091));
    SB_LUT4 Q_15__I_0_add_571_14_lut (.I0(GND_net), .I1(n843_adj_1991[11]), 
            .I2(n668_adj_1716), .I3(n16089), .O(n842_adj_1990[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_14 (.CI(n16089), .I0(n843_adj_1991[11]), 
            .I1(n668_adj_1716), .CO(n16090));
    SB_LUT4 Q_15__I_0_add_571_13_lut (.I0(GND_net), .I1(n843_adj_1991[10]), 
            .I2(n619_adj_268), .I3(n16088), .O(n842_adj_1990[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_13 (.CI(n16088), .I0(n843_adj_1991[10]), 
            .I1(n619_adj_268), .CO(n16089));
    SB_LUT4 Q_15__I_0_add_571_12_lut (.I0(GND_net), .I1(n843_adj_1991[9]), 
            .I2(n570), .I3(n16087), .O(n842_adj_1990[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_12 (.CI(n16087), .I0(n843_adj_1991[9]), .I1(n570), 
            .CO(n16088));
    SB_LUT4 Q_15__I_0_add_571_11_lut (.I0(GND_net), .I1(n843_adj_1991[8]), 
            .I2(n521_adj_1722), .I3(n16086), .O(n842_adj_1990[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_11 (.CI(n16086), .I0(n843_adj_1991[8]), .I1(n521_adj_1722), 
            .CO(n16087));
    SB_LUT4 Q_15__I_0_add_571_10_lut (.I0(GND_net), .I1(n843_adj_1991[7]), 
            .I2(n472_adj_1724), .I3(n16085), .O(n842_adj_1990[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_10 (.CI(n16085), .I0(n843_adj_1991[7]), .I1(n472_adj_1724), 
            .CO(n16086));
    SB_LUT4 Q_15__I_0_add_571_9_lut (.I0(GND_net), .I1(n843_adj_1991[6]), 
            .I2(n423_adj_269), .I3(n16084), .O(n842_adj_1990[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_9 (.CI(n16084), .I0(n843_adj_1991[6]), .I1(n423_adj_269), 
            .CO(n16085));
    SB_LUT4 Q_15__I_0_add_571_8_lut (.I0(GND_net), .I1(n843_adj_1991[5]), 
            .I2(n374_adj_1728), .I3(n16083), .O(n842_adj_1990[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_8 (.CI(n16083), .I0(n843_adj_1991[5]), .I1(n374_adj_1728), 
            .CO(n16084));
    SB_LUT4 Q_15__I_0_add_571_7_lut (.I0(GND_net), .I1(n843_adj_1991[4]), 
            .I2(n325_adj_1730), .I3(n16082), .O(n842_adj_1990[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_7 (.CI(n16082), .I0(n843_adj_1991[4]), .I1(n325_adj_1730), 
            .CO(n16083));
    SB_LUT4 Q_15__I_0_add_571_6_lut (.I0(GND_net), .I1(n843_adj_1991[3]), 
            .I2(n276_adj_270), .I3(n16081), .O(n842_adj_1990[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_6 (.CI(n16081), .I0(n843_adj_1991[3]), .I1(n276_adj_270), 
            .CO(n16082));
    SB_LUT4 Q_15__I_0_add_571_5_lut (.I0(GND_net), .I1(n843_adj_1991[2]), 
            .I2(n227_adj_1734), .I3(n16080), .O(n842_adj_1990[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_5 (.CI(n16080), .I0(n843_adj_1991[2]), .I1(n227_adj_1734), 
            .CO(n16081));
    SB_LUT4 Q_15__I_0_add_571_4_lut (.I0(GND_net), .I1(n843_adj_1991[1]), 
            .I2(n178_adj_1736), .I3(n16079), .O(n842_adj_1990[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_4 (.CI(n16079), .I0(n843_adj_1991[1]), .I1(n178_adj_1736), 
            .CO(n16080));
    SB_LUT4 Q_15__I_0_add_571_3_lut (.I0(GND_net), .I1(n843_adj_1991[0]), 
            .I2(n129_adj_271), .I3(n16078), .O(n842_adj_1990[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_3 (.CI(n16078), .I0(n843_adj_1991[0]), .I1(n129_adj_271), 
            .CO(n16079));
    SB_LUT4 Q_15__I_0_add_571_2_lut (.I0(GND_net), .I1(n35_adj_272), .I2(n80_adj_273), 
            .I3(GND_net), .O(n842_adj_1990[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_571_2 (.CI(GND_net), .I0(n35_adj_272), .I1(n80_adj_273), 
            .CO(n16078));
    SB_LUT4 Q_15__I_0_add_572_16_lut (.I0(GND_net), .I1(n844_adj_1992[13]), 
            .I2(n781_adj_274), .I3(n16076), .O(n843_adj_1991[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_16 (.CI(n16076), .I0(n844_adj_1992[13]), 
            .I1(n781_adj_274), .CO(n783_adj_1744));
    SB_LUT4 Q_15__I_0_add_572_15_lut (.I0(GND_net), .I1(n844_adj_1992[12]), 
            .I2(n720_adj_1746), .I3(n16075), .O(n843_adj_1991[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_15 (.CI(n16075), .I0(n844_adj_1992[12]), 
            .I1(n720_adj_1746), .CO(n16076));
    SB_LUT4 Q_15__I_0_add_572_14_lut (.I0(GND_net), .I1(n844_adj_1992[11]), 
            .I2(n671_adj_1748), .I3(n16074), .O(n843_adj_1991[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_9 (.CI(n16876), .I0(n834[6]), .I1(n396_adj_257), 
            .CO(n16877));
    SB_CARRY Q_15__I_0_add_572_14 (.CI(n16074), .I0(n844_adj_1992[11]), 
            .I1(n671_adj_1748), .CO(n16075));
    SB_LUT4 Q_15__I_0_add_572_13_lut (.I0(GND_net), .I1(n844_adj_1992[10]), 
            .I2(n622_adj_275), .I3(n16073), .O(n843_adj_1991[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_13 (.CI(n16073), .I0(n844_adj_1992[10]), 
            .I1(n622_adj_275), .CO(n16074));
    SB_LUT4 D_15__I_0_10_add_562_8_lut (.I0(GND_net), .I1(n834[5]), .I2(n347_adj_1751), 
            .I3(n16875), .O(n833[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_4 (.CI(n16886), .I0(n833[1]), .I1(n148_adj_1673), 
            .CO(n16887));
    SB_LUT4 Q_15__I_0_add_572_12_lut (.I0(GND_net), .I1(n844_adj_1992[9]), 
            .I2(n573), .I3(n16072), .O(n843_adj_1991[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_12 (.CI(n16072), .I0(n844_adj_1992[9]), .I1(n573), 
            .CO(n16073));
    SB_LUT4 Q_15__I_0_add_572_11_lut (.I0(GND_net), .I1(n844_adj_1992[8]), 
            .I2(n524_adj_1755), .I3(n16071), .O(n843_adj_1991[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_11 (.CI(n16071), .I0(n844_adj_1992[8]), .I1(n524_adj_1755), 
            .CO(n16072));
    SB_LUT4 Q_15__I_0_add_572_10_lut (.I0(GND_net), .I1(n844_adj_1992[7]), 
            .I2(n475_adj_1757), .I3(n16070), .O(n843_adj_1991[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_10 (.CI(n16070), .I0(n844_adj_1992[7]), .I1(n475_adj_1757), 
            .CO(n16071));
    SB_LUT4 Q_15__I_0_add_572_9_lut (.I0(GND_net), .I1(n844_adj_1992[6]), 
            .I2(n426), .I3(n16069), .O(n843_adj_1991[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_9 (.CI(n16069), .I0(n844_adj_1992[6]), .I1(n426), 
            .CO(n16070));
    SB_LUT4 Q_15__I_0_add_572_8_lut (.I0(GND_net), .I1(n844_adj_1992[5]), 
            .I2(n377), .I3(n16068), .O(n843_adj_1991[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_8 (.CI(n16068), .I0(n844_adj_1992[5]), .I1(n377), 
            .CO(n16069));
    SB_LUT4 Q_15__I_0_add_572_7_lut (.I0(GND_net), .I1(n844_adj_1992[4]), 
            .I2(n328), .I3(n16067), .O(n843_adj_1991[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_7 (.CI(n16067), .I0(n844_adj_1992[4]), .I1(n328), 
            .CO(n16068));
    SB_LUT4 Q_15__I_0_add_572_6_lut (.I0(GND_net), .I1(n844_adj_1992[3]), 
            .I2(n279), .I3(n16066), .O(n843_adj_1991[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_6 (.CI(n16066), .I0(n844_adj_1992[3]), .I1(n279), 
            .CO(n16067));
    SB_LUT4 Q_15__I_0_add_572_5_lut (.I0(GND_net), .I1(n844_adj_1992[2]), 
            .I2(n230_c), .I3(n16065), .O(n843_adj_1991[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_5 (.CI(n16065), .I0(n844_adj_1992[2]), .I1(n230_c), 
            .CO(n16066));
    SB_LUT4 Q_15__I_0_add_572_4_lut (.I0(GND_net), .I1(n844_adj_1992[1]), 
            .I2(n181), .I3(n16064), .O(n843_adj_1991[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_4 (.CI(n16064), .I0(n844_adj_1992[1]), .I1(n181), 
            .CO(n16065));
    SB_LUT4 Q_15__I_0_add_572_3_lut (.I0(GND_net), .I1(n844_adj_1992[0]), 
            .I2(n132), .I3(n16063), .O(n843_adj_1991[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_3 (.CI(n16063), .I0(n844_adj_1992[0]), .I1(n132), 
            .CO(n16064));
    SB_LUT4 Q_15__I_0_add_572_2_lut (.I0(GND_net), .I1(n38), .I2(n83), 
            .I3(GND_net), .O(n843_adj_1991[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_572_2 (.CI(GND_net), .I0(n38), .I1(n83), .CO(n16063));
    SB_LUT4 Q_15__I_0_add_573_16_lut (.I0(GND_net), .I1(n845_adj_1993[13]), 
            .I2(n785), .I3(n16061), .O(n844_adj_1992[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_16 (.CI(n16061), .I0(n845_adj_1993[13]), 
            .I1(n785), .CO(n787_adj_1767));
    SB_LUT4 Q_15__I_0_add_573_15_lut (.I0(GND_net), .I1(n845_adj_1993[12]), 
            .I2(n723_adj_1769), .I3(n16060), .O(n844_adj_1992[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_15 (.CI(n16060), .I0(n845_adj_1993[12]), 
            .I1(n723_adj_1769), .CO(n16061));
    SB_LUT4 Q_15__I_0_add_573_14_lut (.I0(GND_net), .I1(n845_adj_1993[11]), 
            .I2(n674_adj_1771), .I3(n16059), .O(n844_adj_1992[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_14 (.CI(n16059), .I0(n845_adj_1993[11]), 
            .I1(n674_adj_1771), .CO(n16060));
    SB_LUT4 Q_15__I_0_add_573_13_lut (.I0(GND_net), .I1(n845_adj_1993[10]), 
            .I2(n625), .I3(n16058), .O(n844_adj_1992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_13 (.CI(n16058), .I0(n845_adj_1993[10]), 
            .I1(n625), .CO(n16059));
    SB_LUT4 Q_15__I_0_add_573_12_lut (.I0(GND_net), .I1(n845_adj_1993[9]), 
            .I2(n576_adj_276), .I3(n16057), .O(n844_adj_1992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_13_lut (.I0(GND_net), .I1(n833[10]), .I2(n589_adj_277), 
            .I3(n16895), .O(Product1_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_12 (.CI(n16057), .I0(n845_adj_1993[9]), .I1(n576_adj_276), 
            .CO(n16058));
    SB_LUT4 Q_15__I_0_add_573_11_lut (.I0(GND_net), .I1(n845_adj_1993[8]), 
            .I2(n527_adj_1778), .I3(n16056), .O(n844_adj_1992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_11 (.CI(n16056), .I0(n845_adj_1993[8]), .I1(n527_adj_1778), 
            .CO(n16057));
    SB_LUT4 Q_15__I_0_add_573_10_lut (.I0(GND_net), .I1(n845_adj_1993[7]), 
            .I2(n478_adj_1780), .I3(n16055), .O(n844_adj_1992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_10 (.CI(n16055), .I0(n845_adj_1993[7]), .I1(n478_adj_1780), 
            .CO(n16056));
    SB_LUT4 Q_15__I_0_add_573_9_lut (.I0(GND_net), .I1(n845_adj_1993[6]), 
            .I2(n429), .I3(n16054), .O(n844_adj_1992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_9 (.CI(n16054), .I0(n845_adj_1993[6]), .I1(n429), 
            .CO(n16055));
    SB_LUT4 Q_15__I_0_add_573_8_lut (.I0(GND_net), .I1(n845_adj_1993[5]), 
            .I2(n380_adj_1784), .I3(n16053), .O(n844_adj_1992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_8 (.CI(n16053), .I0(n845_adj_1993[5]), .I1(n380_adj_1784), 
            .CO(n16054));
    SB_LUT4 Q_15__I_0_add_573_7_lut (.I0(GND_net), .I1(n845_adj_1993[4]), 
            .I2(n331_adj_1786), .I3(n16052), .O(n844_adj_1992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_7 (.CI(n16052), .I0(n845_adj_1993[4]), .I1(n331_adj_1786), 
            .CO(n16053));
    SB_LUT4 Q_15__I_0_add_573_6_lut (.I0(GND_net), .I1(n845_adj_1993[3]), 
            .I2(n282), .I3(n16051), .O(n844_adj_1992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_6 (.CI(n16051), .I0(n845_adj_1993[3]), .I1(n282), 
            .CO(n16052));
    SB_LUT4 Q_15__I_0_add_573_5_lut (.I0(GND_net), .I1(n845_adj_1993[2]), 
            .I2(n233_adj_1790), .I3(n16050), .O(n844_adj_1992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_5 (.CI(n16050), .I0(n845_adj_1993[2]), .I1(n233_adj_1790), 
            .CO(n16051));
    SB_LUT4 Q_15__I_0_add_573_4_lut (.I0(GND_net), .I1(n845_adj_1993[1]), 
            .I2(n184_adj_1792), .I3(n16049), .O(n844_adj_1992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_4 (.CI(n16049), .I0(n845_adj_1993[1]), .I1(n184_adj_1792), 
            .CO(n16050));
    SB_LUT4 Q_15__I_0_add_573_3_lut (.I0(GND_net), .I1(n845_adj_1993[0]), 
            .I2(n135), .I3(n16048), .O(n844_adj_1992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_3 (.CI(n16048), .I0(n845_adj_1993[0]), .I1(n135), 
            .CO(n16049));
    SB_LUT4 Q_15__I_0_add_573_2_lut (.I0(GND_net), .I1(n41), .I2(n86_adj_278), 
            .I3(GND_net), .O(n844_adj_1992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_573_2 (.CI(GND_net), .I0(n41), .I1(n86_adj_278), 
            .CO(n16048));
    SB_LUT4 Q_15__I_0_add_574_16_lut (.I0(GND_net), .I1(n846_adj_1994[13]), 
            .I2(n789), .I3(n16046), .O(n845_adj_1993[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_16 (.CI(n16046), .I0(n846_adj_1994[13]), 
            .I1(n789), .CO(n791_adj_1798));
    SB_LUT4 Q_15__I_0_add_574_15_lut (.I0(GND_net), .I1(n846_adj_1994[12]), 
            .I2(n726), .I3(n16045), .O(n845_adj_1993[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_15 (.CI(n16045), .I0(n846_adj_1994[12]), 
            .I1(n726), .CO(n16046));
    SB_LUT4 Q_15__I_0_add_574_14_lut (.I0(GND_net), .I1(n846_adj_1994[11]), 
            .I2(n677), .I3(n16044), .O(n845_adj_1993[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_14 (.CI(n16044), .I0(n846_adj_1994[11]), 
            .I1(n677), .CO(n16045));
    SB_LUT4 Q_15__I_0_add_574_13_lut (.I0(GND_net), .I1(n846_adj_1994[10]), 
            .I2(n628), .I3(n16043), .O(n845_adj_1993[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_13 (.CI(n16043), .I0(n846_adj_1994[10]), 
            .I1(n628), .CO(n16044));
    SB_LUT4 Q_15__I_0_add_574_12_lut (.I0(GND_net), .I1(n846_adj_1994[9]), 
            .I2(n579), .I3(n16042), .O(n845_adj_1993[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_12 (.CI(n16042), .I0(n846_adj_1994[9]), .I1(n579), 
            .CO(n16043));
    SB_LUT4 Q_15__I_0_add_574_11_lut (.I0(GND_net), .I1(n846_adj_1994[8]), 
            .I2(n530), .I3(n16041), .O(n845_adj_1993[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_11 (.CI(n16041), .I0(n846_adj_1994[8]), .I1(n530), 
            .CO(n16042));
    SB_LUT4 Q_15__I_0_add_574_10_lut (.I0(GND_net), .I1(n846_adj_1994[7]), 
            .I2(n481), .I3(n16040), .O(n845_adj_1993[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_10 (.CI(n16040), .I0(n846_adj_1994[7]), .I1(n481), 
            .CO(n16041));
    SB_LUT4 Q_15__I_0_add_574_9_lut (.I0(GND_net), .I1(n846_adj_1994[6]), 
            .I2(n432), .I3(n16039), .O(n845_adj_1993[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_9 (.CI(n16039), .I0(n846_adj_1994[6]), .I1(n432), 
            .CO(n16040));
    SB_LUT4 Q_15__I_0_add_574_8_lut (.I0(GND_net), .I1(n846_adj_1994[5]), 
            .I2(n383), .I3(n16038), .O(n845_adj_1993[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_8 (.CI(n16038), .I0(n846_adj_1994[5]), .I1(n383), 
            .CO(n16039));
    SB_LUT4 Q_15__I_0_add_574_7_lut (.I0(GND_net), .I1(n846_adj_1994[4]), 
            .I2(n334), .I3(n16037), .O(n845_adj_1993[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_7 (.CI(n16037), .I0(n846_adj_1994[4]), .I1(n334), 
            .CO(n16038));
    SB_LUT4 Q_15__I_0_add_574_6_lut (.I0(GND_net), .I1(n846_adj_1994[3]), 
            .I2(n285), .I3(n16036), .O(n845_adj_1993[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_6 (.CI(n16036), .I0(n846_adj_1994[3]), .I1(n285), 
            .CO(n16037));
    SB_LUT4 Q_15__I_0_add_574_5_lut (.I0(GND_net), .I1(n846_adj_1994[2]), 
            .I2(n236_adj_1810), .I3(n16035), .O(n845_adj_1993[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_5 (.CI(n16035), .I0(n846_adj_1994[2]), .I1(n236_adj_1810), 
            .CO(n16036));
    SB_LUT4 Q_15__I_0_add_574_4_lut (.I0(GND_net), .I1(n846_adj_1994[1]), 
            .I2(n187_adj_1812), .I3(n16034), .O(n845_adj_1993[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_4 (.CI(n16034), .I0(n846_adj_1994[1]), .I1(n187_adj_1812), 
            .CO(n16035));
    SB_LUT4 Q_15__I_0_add_574_3_lut (.I0(GND_net), .I1(n846_adj_1994[0]), 
            .I2(n138_adj_279), .I3(n16033), .O(n845_adj_1993[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_3 (.CI(n16033), .I0(n846_adj_1994[0]), .I1(n138_adj_279), 
            .CO(n16034));
    SB_LUT4 Q_15__I_0_add_574_2_lut (.I0(GND_net), .I1(n44_adj_280), .I2(n89_adj_281), 
            .I3(GND_net), .O(n845_adj_1993[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_574_2 (.CI(GND_net), .I0(n44_adj_280), .I1(n89_adj_281), 
            .CO(n16033));
    SB_LUT4 Q_15__I_0_add_575_16_lut (.I0(GND_net), .I1(n19580), .I2(n19604), 
            .I3(n16032), .O(n846_adj_1994[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_add_575_15_lut (.I0(GND_net), .I1(n685_adj_282), .I2(n729_adj_1819), 
            .I3(n16031), .O(n846_adj_1994[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_15 (.CI(n16031), .I0(n685_adj_282), .I1(n729_adj_1819), 
            .CO(n16032));
    SB_LUT4 Q_15__I_0_add_575_14_lut (.I0(GND_net), .I1(n636_adj_1820), 
            .I2(n680_adj_1821), .I3(n16030), .O(n846_adj_1994[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_14 (.CI(n16030), .I0(n636_adj_1820), .I1(n680_adj_1821), 
            .CO(n16031));
    SB_LUT4 Q_15__I_0_add_575_13_lut (.I0(GND_net), .I1(n587_adj_283), .I2(n631_adj_284), 
            .I3(n16029), .O(n846_adj_1994[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_13 (.CI(n16029), .I0(n587_adj_283), .I1(n631_adj_284), 
            .CO(n16030));
    SB_LUT4 Q_15__I_0_add_575_12_lut (.I0(GND_net), .I1(n538_adj_285), .I2(n582), 
            .I3(n16028), .O(n846_adj_1994[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_12 (.CI(n16028), .I0(n538_adj_285), .I1(n582), 
            .CO(n16029));
    SB_LUT4 Q_15__I_0_add_575_11_lut (.I0(GND_net), .I1(n489_adj_286), .I2(n533_adj_1827), 
            .I3(n16027), .O(n846_adj_1994[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_11 (.CI(n16027), .I0(n489_adj_286), .I1(n533_adj_1827), 
            .CO(n16028));
    SB_LUT4 Q_15__I_0_add_575_10_lut (.I0(GND_net), .I1(n440_adj_1828), 
            .I2(n484_adj_1829), .I3(n16026), .O(n846_adj_1994[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_10 (.CI(n16026), .I0(n440_adj_1828), .I1(n484_adj_1829), 
            .CO(n16027));
    SB_LUT4 Q_15__I_0_add_575_9_lut (.I0(GND_net), .I1(n391_adj_287), .I2(n435_adj_288), 
            .I3(n16025), .O(n846_adj_1994[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_9 (.CI(n16025), .I0(n391_adj_287), .I1(n435_adj_288), 
            .CO(n16026));
    SB_LUT4 Q_15__I_0_add_575_8_lut (.I0(GND_net), .I1(n342_adj_289), .I2(n386_adj_1833), 
            .I3(n16024), .O(n846_adj_1994[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_8 (.CI(n16024), .I0(n342_adj_289), .I1(n386_adj_1833), 
            .CO(n16025));
    SB_LUT4 Q_15__I_0_add_575_7_lut (.I0(GND_net), .I1(n293_adj_1834), .I2(n337_adj_1835), 
            .I3(n16023), .O(n846_adj_1994[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_7 (.CI(n16023), .I0(n293_adj_1834), .I1(n337_adj_1835), 
            .CO(n16024));
    SB_LUT4 Q_15__I_0_add_575_6_lut (.I0(GND_net), .I1(n244_adj_290), .I2(n288_adj_291), 
            .I3(n16022), .O(n846_adj_1994[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_6 (.CI(n16022), .I0(n244_adj_290), .I1(n288_adj_291), 
            .CO(n16023));
    SB_LUT4 Q_15__I_0_add_575_5_lut (.I0(GND_net), .I1(n195_adj_292), .I2(n239_adj_1839), 
            .I3(n16021), .O(n846_adj_1994[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_5 (.CI(n16021), .I0(n195_adj_292), .I1(n239_adj_1839), 
            .CO(n16022));
    SB_LUT4 Q_15__I_0_add_575_4_lut (.I0(GND_net), .I1(n146_adj_1840), .I2(n190_adj_1841), 
            .I3(n16020), .O(n846_adj_1994[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_4 (.CI(n16020), .I0(n146_adj_1840), .I1(n190_adj_1841), 
            .CO(n16021));
    SB_LUT4 Q_15__I_0_add_575_3_lut (.I0(GND_net), .I1(n97_adj_1842), .I2(n141_adj_293), 
            .I3(n16019), .O(n846_adj_1994[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_3 (.CI(n16019), .I0(n97_adj_1842), .I1(n141_adj_293), 
            .CO(n16020));
    SB_LUT4 Q_15__I_0_add_575_2_lut (.I0(GND_net), .I1(n48_adj_1844), .I2(n92_adj_294), 
            .I3(GND_net), .O(n846_adj_1994[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_add_575_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_add_575_2 (.CI(GND_net), .I0(n48_adj_1844), .I1(n92_adj_294), 
            .CO(n16019));
    SB_LUT4 add_1227_16_lut (.I0(GND_net), .I1(n846_adj_1994[14]), .I2(n791_adj_1798), 
            .I3(n16018), .O(Product4_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1227_15_lut (.I0(GND_net), .I1(n845_adj_1993[14]), .I2(n787_adj_1767), 
            .I3(n16017), .O(Product4_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_15 (.CI(n16017), .I0(n845_adj_1993[14]), .I1(n787_adj_1767), 
            .CO(n16018));
    SB_LUT4 add_1227_14_lut (.I0(GND_net), .I1(n844_adj_1992[14]), .I2(n783_adj_1744), 
            .I3(n16016), .O(Product4_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_14 (.CI(n16016), .I0(n844_adj_1992[14]), .I1(n783_adj_1744), 
            .CO(n16017));
    SB_LUT4 add_1227_13_lut (.I0(GND_net), .I1(n843_adj_1991[14]), .I2(n779_adj_1712), 
            .I3(n16015), .O(Product4_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_13 (.CI(n16015), .I0(n843_adj_1991[14]), .I1(n779_adj_1712), 
            .CO(n16016));
    SB_LUT4 add_1227_12_lut (.I0(GND_net), .I1(n842_adj_1990[14]), .I2(n775_adj_1680), 
            .I3(n16014), .O(Product4_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_12 (.CI(n16014), .I0(n842_adj_1990[14]), .I1(n775_adj_1680), 
            .CO(n16015));
    SB_LUT4 add_1227_11_lut (.I0(GND_net), .I1(n841_adj_1989[14]), .I2(n771_adj_1561), 
            .I3(n16013), .O(Product4_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_11 (.CI(n16013), .I0(n841_adj_1989[14]), .I1(n771_adj_1561), 
            .CO(n16014));
    SB_LUT4 add_1227_10_lut (.I0(GND_net), .I1(n840_adj_1988[14]), .I2(n767_adj_1523), 
            .I3(n16012), .O(Product4_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_10 (.CI(n16012), .I0(n840_adj_1988[14]), .I1(n767_adj_1523), 
            .CO(n16013));
    SB_LUT4 add_1227_9_lut (.I0(GND_net), .I1(n839_adj_1987[14]), .I2(n763_adj_1502), 
            .I3(n16011), .O(Product4_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_9 (.CI(n16011), .I0(n839_adj_1987[14]), .I1(n763_adj_1502), 
            .CO(n16012));
    SB_LUT4 add_1227_8_lut (.I0(GND_net), .I1(n838_adj_1986[14]), .I2(n759_adj_1482), 
            .I3(n16010), .O(Product4_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_8 (.CI(n16010), .I0(n838_adj_1986[14]), .I1(n759_adj_1482), 
            .CO(n16011));
    SB_LUT4 add_1227_7_lut (.I0(GND_net), .I1(n837_adj_1985[14]), .I2(n755_adj_1464), 
            .I3(n16009), .O(Product4_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_7 (.CI(n16009), .I0(n837_adj_1985[14]), .I1(n755_adj_1464), 
            .CO(n16010));
    SB_LUT4 add_1227_6_lut (.I0(GND_net), .I1(n836_adj_1984[14]), .I2(n751_adj_1446), 
            .I3(n16008), .O(Product4_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_6 (.CI(n16008), .I0(n836_adj_1984[14]), .I1(n751_adj_1446), 
            .CO(n16009));
    SB_LUT4 add_1227_5_lut (.I0(GND_net), .I1(n835_adj_1983[14]), .I2(n747_adj_1425), 
            .I3(n16007), .O(Product4_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_5 (.CI(n16007), .I0(n835_adj_1983[14]), .I1(n747_adj_1425), 
            .CO(n16008));
    SB_LUT4 add_1227_4_lut (.I0(GND_net), .I1(n834_adj_1982[14]), .I2(n743_adj_1411), 
            .I3(n16006), .O(Product4_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_4 (.CI(n16006), .I0(n834_adj_1982[14]), .I1(n743_adj_1411), 
            .CO(n16007));
    SB_LUT4 add_1227_3_lut (.I0(GND_net), .I1(n833_adj_1981[14]), .I2(n739_adj_1396), 
            .I3(n16005), .O(Product4_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_3 (.CI(n16005), .I0(n833_adj_1981[14]), .I1(n739_adj_1396), 
            .CO(n16006));
    SB_LUT4 add_1227_2_lut (.I0(GND_net), .I1(\qVoltage[15] ), .I2(Look_Up_Table_out1_1[15]), 
            .I3(n16004), .O(Product4_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1227_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1227_2 (.CI(n16004), .I0(\qVoltage[15] ), .I1(Look_Up_Table_out1_1[15]), 
            .CO(n16005));
    SB_CARRY add_1227_1 (.CI(GND_net), .I0(n832_adj_1980[14]), .I1(n832_adj_1980[14]), 
            .CO(n16004));
    SB_LUT4 add_7655_25_lut (.I0(GND_net), .I1(Product3_mul_temp[25]), .I2(Product4_mul_temp[25]), 
            .I3(n17691), .O(\betaVoltage[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_7 (.CI(n16560), .I0(n842[4]), .I1(n331), 
            .CO(n16561));
    SB_CARRY Q_15__I_0_11_add_563_16 (.CI(n16674), .I0(n835[13]), .I1(n793), 
            .CO(n747_adj_1337));
    SB_CARRY add_7655_25 (.CI(n17691), .I0(Product3_mul_temp[25]), .I1(Product4_mul_temp[25]), 
            .CO(n17692));
    SB_LUT4 Q_15__I_0_11_add_570_6_lut (.I0(GND_net), .I1(n842[3]), .I2(n282_c), 
            .I3(n16559), .O(n841_adj_1952[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_15_lut (.I0(GND_net), .I1(n835[12]), .I2(n723), 
            .I3(n16673), .O(n834_adj_1976[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_6 (.CI(n16559), .I0(n842[3]), .I1(n282_c), 
            .CO(n16560));
    SB_LUT4 D_15__I_0_10_i377_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n558_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7336_2_lut (.I0(n833_adj_1964[13]), .I1(\dVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n9108));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam i7336_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7756_2_lut (.I0(n834_adj_1962[13]), .I1(\dVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n833_adj_1964[14]));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam i7756_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7758_2_lut (.I0(n834_adj_1962[13]), .I1(\dVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n9531));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam i7758_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_563_6 (.CI(n16858), .I0(n835_adj_1961[3]), 
            .I1(n252_adj_256), .CO(n16859));
    SB_LUT4 D_15__I_0_10_add_563_5_lut (.I0(GND_net), .I1(n835_adj_1961[2]), 
            .I2(n203), .I3(n16857), .O(n834[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_14_lut (.I0(GND_net), .I1(n835_adj_1961[11]), 
            .I2(n644_adj_1851), .I3(n16866), .O(n834[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_8 (.CI(n16875), .I0(n834[5]), .I1(n347_adj_1751), 
            .CO(n16876));
    SB_LUT4 D_15__I_0_10_add_561_3_lut (.I0(GND_net), .I1(n833[0]), .I2(n99_adj_295), 
            .I3(n16885), .O(Product1_mul_temp[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_3 (.CI(n16885), .I0(n833[0]), .I1(n99_adj_295), 
            .CO(n16886));
    SB_LUT4 D_15__I_0_10_i470_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n696_adj_1380));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i470_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i233_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_1377));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i261_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n386));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i367_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n543_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i303_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_1374));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i303_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_561_13 (.CI(n16895), .I0(n833[10]), .I1(n589_adj_277), 
            .CO(n16896));
    SB_LUT4 D_15__I_0_10_i387_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n573_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i387_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i113_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n166));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i342_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n506_adj_1370));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i342_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i439_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n650_adj_1366));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i439_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i472_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n699_adj_1363));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i472_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i307_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_1361));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i307_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i109_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n160_adj_1359));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i375_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n555_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_566_7 (.CI(n16814), .I0(n838[4]), .I1(n310_adj_1660), 
            .CO(n16815));
    SB_LUT4 D_15__I_0_10_i255_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n377_adj_1853));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_567_2 (.CI(GND_net), .I0(n23_adj_254), .I1(n68_adj_255), 
            .CO(n16795));
    SB_LUT4 D_15__I_0_10_add_564_12_lut (.I0(GND_net), .I1(n836_adj_1960[9]), 
            .I2(n549_adj_1662), .I3(n16849), .O(n835_adj_1961[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_13 (.CI(n16850), .I0(n836_adj_1960[10]), 
            .I1(n598), .CO(n16851));
    SB_LUT4 add_7655_24_lut (.I0(GND_net), .I1(Product3_mul_temp[24]), .I2(Product4_mul_temp[24]), 
            .I3(n17690), .O(\betaVoltage[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_563_5 (.CI(n16857), .I0(n835_adj_1961[2]), 
            .I1(n203), .CO(n16858));
    SB_LUT4 D_15__I_0_10_i474_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n702_adj_1855));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i474_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_563_14 (.CI(n16866), .I0(n835_adj_1961[11]), 
            .I1(n644_adj_1851), .CO(n16867));
    SB_LUT4 D_15__I_0_10_add_562_7_lut (.I0(GND_net), .I1(n834[4]), .I2(n298_adj_1856), 
            .I3(n16874), .O(n833[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_7 (.CI(n16874), .I0(n834[4]), .I1(n298_adj_1856), 
            .CO(n16875));
    SB_CARRY Q_15__I_0_11_add_563_15 (.CI(n16673), .I0(n835[12]), .I1(n723), 
            .CO(n16674));
    SB_LUT4 Q_15__I_0_11_add_570_5_lut (.I0(GND_net), .I1(n842[2]), .I2(n233_c), 
            .I3(n16558), .O(n841_adj_1952[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_14_lut (.I0(GND_net), .I1(n835[11]), .I2(n674), 
            .I3(n16672), .O(n833_adj_1977[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_24 (.CI(n17690), .I0(Product3_mul_temp[24]), .I1(Product4_mul_temp[24]), 
            .CO(n17691));
    SB_LUT4 D_15__I_0_10_i433_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n641_adj_1353));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i433_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_561_2 (.CI(GND_net), .I0(n19576), .I1(n50_adj_296), 
            .CO(n16885));
    SB_LUT4 add_7655_23_lut (.I0(GND_net), .I1(Product3_mul_temp[23]), .I2(Product4_mul_temp[23]), 
            .I3(n17689), .O(\betaVoltage[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_561_12_lut (.I0(GND_net), .I1(n833[9]), .I2(n540_adj_1860), 
            .I3(n16894), .O(Product1_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_10 (.CI(n16593), .I0(n840[7]), .I1(n478), 
            .CO(n16594));
    SB_CARRY add_7655_23 (.CI(n17689), .I0(Product3_mul_temp[23]), .I1(Product4_mul_temp[23]), 
            .CO(n17690));
    SB_CARRY Q_15__I_0_11_add_563_14 (.CI(n16672), .I0(n835[11]), .I1(n674), 
            .CO(n16673));
    SB_LUT4 Q_15__I_0_11_add_568_9_lut (.I0(GND_net), .I1(n840[6]), .I2(n429_c), 
            .I3(n16592), .O(n839[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_13_lut (.I0(GND_net), .I1(n835[10]), .I2(n625_c), 
            .I3(n16671), .O(Product2_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_570_5 (.CI(n16558), .I0(n842[2]), .I1(n233_c), 
            .CO(n16559));
    SB_LUT4 D_15__I_0_10_i105_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n154_adj_1862));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i365_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n540_adj_1860));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7439_2_lut (.I0(n833_adj_1977[13]), .I1(\qVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n832_adj_1978[14]));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam i7439_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 D_15__I_0_10_i336_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n497_adj_1351));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i336_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i202_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n298_adj_1856));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_add_566_6_lut (.I0(GND_net), .I1(n838[3]), .I2(n261_adj_297), 
            .I3(n16813), .O(n837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_14 (.CI(n16806), .I0(n839_adj_1951[11]), 
            .I1(n656_adj_1646), .CO(n16807));
    SB_CARRY D_15__I_0_10_add_572_10 (.CI(n16727), .I0(n844_adj_1959[7]), 
            .I1(n475), .CO(n16728));
    SB_LUT4 D_15__I_0_10_i435_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n644_adj_1851));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i435_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i445_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n659));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i33_2_lut (.I0(n19702), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n48_adj_1844));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i33_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_add_563_4_lut (.I0(GND_net), .I1(n835_adj_1961[1]), 
            .I2(n154_adj_1862), .I3(n16856), .O(n834[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_13_lut (.I0(GND_net), .I1(n835_adj_1961[10]), 
            .I2(n595_adj_298), .I3(n16865), .O(n834[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_562_6_lut (.I0(GND_net), .I1(n834[3]), .I2(n249_adj_299), 
            .I3(n16873), .O(n833[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_6 (.CI(n16873), .I0(n834[3]), .I1(n249_adj_299), 
            .CO(n16874));
    SB_LUT4 D_15__I_0_10_add_562_16_lut (.I0(GND_net), .I1(n834[13]), .I2(n741_adj_300), 
            .I3(n16883), .O(n833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_12 (.CI(n16894), .I0(n833[9]), .I1(n540_adj_1860), 
            .CO(n16895));
    SB_LUT4 i3_4_lut (.I0(Out_31__N_333), .I1(\preSatVoltage[10] ), .I2(Out_31__N_332), 
            .I3(Look_Up_Table_out1_1[15]), .O(n97_adj_1842));
    defparam i3_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i7441_2_lut (.I0(n833_adj_1977[13]), .I1(\qVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n9213));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam i7441_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7861_2_lut (.I0(n834_adj_1976[13]), .I1(\qVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n833_adj_1977[14]));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam i7861_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 Q_15__I_0_i129_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n190_adj_1841));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i129_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i99_2_lut (.I0(\qVoltage[2] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n146_adj_1840));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i99_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_i453_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n671));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i162_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n239_adj_1839));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i228_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n337_adj_1835));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i198_2_lut (.I0(\qVoltage[5] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_1834));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i198_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i7863_2_lut (.I0(n834_adj_1976[13]), .I1(\qVoltage[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n9636));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam i7863_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i261_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n386_adj_1833));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i327_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_1829));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i297_2_lut (.I0(\qVoltage[8] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n440_adj_1828));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i297_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_i360_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_1827));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i360_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i327_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i297_2_lut (.I0(\dVoltage[8] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n440_adj_1341));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i297_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_i360_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i360_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i459_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n680_adj_1821));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i429_2_lut (.I0(\qVoltage[12] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n636_adj_1820));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i429_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_i492_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n729_adj_1819));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i492_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_566_16 (.CI(n16823), .I0(n838[13]), .I1(n757_adj_253), 
            .CO(n759));
    SB_LUT4 D_15__I_0_10_add_566_15_lut (.I0(GND_net), .I1(n838[12]), .I2(n702_adj_1855), 
            .I3(n16822), .O(n837[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_13 (.CI(n16671), .I0(n835[10]), .I1(n625_c), 
            .CO(n16672));
    SB_LUT4 D_15__I_0_10_i486_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n720));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i486_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_565_7 (.CI(n16829), .I0(n837[4]), .I1(n307_adj_1653), 
            .CO(n16830));
    SB_LUT4 Q_15__I_0_11_add_570_4_lut (.I0(GND_net), .I1(n842[1]), .I2(n184), 
            .I3(n16557), .O(n841_adj_1952[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_12_lut (.I0(GND_net), .I1(n835[9]), .I2(n576), 
            .I3(n16670), .O(Product2_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_572_9_lut (.I0(GND_net), .I1(n844_adj_1959[6]), 
            .I2(n426_adj_301), .I3(n16726), .O(n843_adj_1956[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_9 (.CI(n16726), .I0(n844_adj_1959[6]), 
            .I1(n426_adj_301), .CO(n16727));
    SB_CARRY Q_15__I_0_11_add_570_4 (.CI(n16557), .I0(n842[1]), .I1(n184), 
            .CO(n16558));
    SB_LUT4 D_15__I_0_10_add_572_8_lut (.I0(GND_net), .I1(n844_adj_1959[5]), 
            .I2(n377_adj_1853), .I3(n16725), .O(n843_adj_1956[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_12 (.CI(n16670), .I0(n835[9]), .I1(n576), 
            .CO(n16671));
    SB_CARRY Q_15__I_0_11_add_566_13 (.CI(n16626), .I0(n838_adj_1953[10]), 
            .I1(n625_c), .CO(n16627));
    SB_CARRY D_15__I_0_10_add_572_8 (.CI(n16725), .I0(n844_adj_1959[5]), 
            .I1(n377_adj_1853), .CO(n16726));
    SB_LUT4 D_15__I_0_10_add_565_6_lut (.I0(GND_net), .I1(n837[3]), .I2(n258_adj_302), 
            .I3(n16828), .O(n836_adj_1960[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(Out_31__N_332), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[13] ), .O(n244_c));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h4044;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_294 (.I0(Out_31__N_332), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[12] ), .O(n195_c));
    defparam i1_2_lut_3_lut_4_lut_adj_294.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_i127_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n187_adj_1812));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i127_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_295 (.I0(Out_31__N_332), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[19] ), .O(n538_c));
    defparam i1_2_lut_3_lut_4_lut_adj_295.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_i160_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n236_adj_1810));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i127_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n187));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i127_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_296 (.I0(Out_31__N_332), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[22] ), .O(n685_adj_1082));
    defparam i1_2_lut_3_lut_4_lut_adj_296.LUT_INIT = 16'h4044;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_297 (.I0(Out_31__N_332), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[23] ), .O(n19680));
    defparam i1_2_lut_3_lut_4_lut_adj_297.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_i226_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n334));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i259_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n383));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i325_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i325_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i33_2_lut (.I0(n19352), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n48_adj_1326));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i33_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_i358_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i358_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_298 (.I0(Out_31__N_333_adj_303), .I1(\preSatVoltage[10]_adj_304 ), 
            .I2(Out_31__N_332_adj_305), .I3(\Product_mul_temp[26] ), .O(n97_adj_1322));
    defparam i3_4_lut_adj_298.LUT_INIT = 16'h0100;
    SB_LUT4 Q_15__I_0_i457_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n677));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i490_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n726));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i490_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i125_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n184_adj_1792));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i125_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i158_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n233_adj_1790));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i224_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n331_adj_1786));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i257_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n380_adj_1784));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i323_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_1780));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i323_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i99_2_lut (.I0(\dVoltage[2] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n146_adj_1321));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i99_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_i356_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_1778));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i356_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_add_567_9_lut (.I0(GND_net), .I1(n839_adj_1951[6]), 
            .I2(n411_adj_306), .I3(n16801), .O(n838[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_6 (.CI(n16828), .I0(n837[3]), .I1(n258_adj_302), 
            .CO(n16829));
    SB_LUT4 D_15__I_0_10_add_565_11_lut (.I0(GND_net), .I1(n837[8]), .I2(n503_adj_1020), 
            .I3(n16833), .O(n836_adj_1960[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_564_2_lut (.I0(GND_net), .I1(n14_adj_307), 
            .I2(n59_adj_308), .I3(GND_net), .O(n835_adj_1961[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_2 (.CI(GND_net), .I0(n14_adj_307), .I1(n59_adj_308), 
            .CO(n16840));
    SB_CARRY D_15__I_0_10_add_563_4 (.CI(n16856), .I0(n835_adj_1961[1]), 
            .I1(n154_adj_1862), .CO(n16857));
    SB_CARRY D_15__I_0_10_add_563_13 (.CI(n16865), .I0(n835_adj_1961[10]), 
            .I1(n595_adj_298), .CO(n16866));
    SB_LUT4 D_15__I_0_10_add_562_5_lut (.I0(GND_net), .I1(n834[2]), .I2(n200), 
            .I3(n16872), .O(n833[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_5 (.CI(n16872), .I0(n834[2]), .I1(n200), 
            .CO(n16873));
    SB_CARRY D_15__I_0_10_add_564_8 (.CI(n16845), .I0(n836_adj_1960[5]), 
            .I1(n353_adj_1655), .CO(n16846));
    SB_CARRY D_15__I_0_10_add_562_16 (.CI(n16883), .I0(n834[13]), .I1(n741_adj_300), 
            .CO(n743));
    SB_LUT4 D_15__I_0_10_add_561_11_lut (.I0(GND_net), .I1(n833[8]), .I2(n491), 
            .I3(n16893), .O(Product1_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_11 (.CI(n16833), .I0(n837[8]), .I1(n503_adj_1020), 
            .CO(n16834));
    SB_CARRY D_15__I_0_10_add_566_6 (.CI(n16813), .I0(n838[3]), .I1(n261_adj_297), 
            .CO(n16814));
    SB_LUT4 D_15__I_0_10_add_565_16_lut (.I0(GND_net), .I1(n837[13]), .I2(n753_adj_309), 
            .I3(n16838), .O(n836_adj_1960[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_3_lut (.I0(GND_net), .I1(n835_adj_1961[0]), 
            .I2(n105_adj_310), .I3(n16855), .O(n834[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_563_3 (.CI(n16855), .I0(n835_adj_1961[0]), 
            .I1(n105_adj_310), .CO(n16856));
    SB_LUT4 D_15__I_0_10_add_564_7_lut (.I0(GND_net), .I1(n836_adj_1960[4]), 
            .I2(n304), .I3(n16844), .O(n835_adj_1961[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_12_lut (.I0(GND_net), .I1(n835_adj_1961[9]), 
            .I2(n546_c), .I3(n16864), .O(n834[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_564_7 (.CI(n16844), .I0(n836_adj_1960[4]), 
            .I1(n304), .CO(n16845));
    SB_LUT4 D_15__I_0_10_add_562_4_lut (.I0(GND_net), .I1(n834[1]), .I2(n151_adj_1886), 
            .I3(n16871), .O(n833[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_562_15_lut (.I0(GND_net), .I1(n834[12]), .I2(n690_adj_1887), 
            .I3(n16882), .O(n833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_15 (.CI(n16882), .I0(n834[12]), .I1(n690_adj_1887), 
            .CO(n16883));
    SB_LUT4 D_15__I_0_10_add_568_16_lut (.I0(GND_net), .I1(n840_adj_1950[13]), 
            .I2(n765_adj_311), .I3(n16793), .O(n839_adj_1951[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_568_16 (.CI(n16793), .I0(n840_adj_1950[13]), 
            .I1(n765_adj_311), .CO(n767_adj_1092));
    SB_CARRY D_15__I_0_10_add_561_11 (.CI(n16893), .I0(n833[8]), .I1(n491), 
            .CO(n16894));
    SB_LUT4 D_15__I_0_10_add_561_10_lut (.I0(GND_net), .I1(n833[7]), .I2(n442_adj_1889), 
            .I3(n16892), .O(Product1_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_9 (.CI(n16801), .I0(n839_adj_1951[6]), 
            .I1(n411_adj_306), .CO(n16802));
    SB_CARRY D_15__I_0_10_add_566_15 (.CI(n16822), .I0(n838[12]), .I1(n702_adj_1855), 
            .CO(n16823));
    SB_LUT4 D_15__I_0_10_add_566_14_lut (.I0(GND_net), .I1(n838[11]), .I2(n653_adj_1891), 
            .I3(n16821), .O(n837[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_563_2_lut (.I0(GND_net), .I1(n11), .I2(n56), 
            .I3(GND_net), .O(n834[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_563_12 (.CI(n16864), .I0(n835_adj_1961[9]), 
            .I1(n546_c), .CO(n16865));
    SB_LUT4 D_15__I_0_10_add_563_11_lut (.I0(GND_net), .I1(n835_adj_1961[8]), 
            .I2(n497_adj_1351), .I3(n16863), .O(n834[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_562_4 (.CI(n16871), .I0(n834[1]), .I1(n151_adj_1886), 
            .CO(n16872));
    SB_LUT4 D_15__I_0_10_add_562_14_lut (.I0(GND_net), .I1(n834[11]), .I2(n641_adj_1353), 
            .I3(n16881), .O(n833[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_561_10 (.CI(n16892), .I0(n833[7]), .I1(n442_adj_1889), 
            .CO(n16893));
    SB_LUT4 D_15__I_0_10_add_561_9_lut (.I0(GND_net), .I1(n833[6]), .I2(n393), 
            .I3(n16891), .O(Product1_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_8_lut (.I0(GND_net), .I1(n839_adj_1951[5]), 
            .I2(n362_adj_1892), .I3(n16800), .O(n838[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_572_7_lut (.I0(GND_net), .I1(n844_adj_1959[4]), 
            .I2(n328_adj_1894), .I3(n16724), .O(n843_adj_1956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_568_15_lut (.I0(GND_net), .I1(n840_adj_1950[12]), 
            .I2(n708), .I3(n16792), .O(n839_adj_1951[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_567_8 (.CI(n16800), .I0(n839_adj_1951[5]), 
            .I1(n362_adj_1892), .CO(n16801));
    SB_LUT4 D_15__I_0_10_add_567_7_lut (.I0(GND_net), .I1(n839_adj_1951[4]), 
            .I2(n313), .I3(n16799), .O(n838[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_567_13_lut (.I0(GND_net), .I1(n839_adj_1951[10]), 
            .I2(n607_adj_312), .I3(n16805), .O(n838[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_566_5_lut (.I0(GND_net), .I1(n838[2]), .I2(n212), 
            .I3(n16812), .O(n837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_14 (.CI(n16821), .I0(n838[11]), .I1(n653_adj_1891), 
            .CO(n16822));
    SB_LUT4 D_15__I_0_10_add_566_13_lut (.I0(GND_net), .I1(n838[10]), .I2(n604_adj_313), 
            .I3(n16820), .O(n837[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_565_5_lut (.I0(GND_net), .I1(n837[2]), .I2(n209), 
            .I3(n16827), .O(n836_adj_1960[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_565_10_lut (.I0(GND_net), .I1(n837[7]), .I2(n454_adj_1361), 
            .I3(n16832), .O(n836_adj_1960[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_565_16 (.CI(n16838), .I0(n837[13]), .I1(n753_adj_309), 
            .CO(n755_adj_1094));
    SB_LUT4 D_15__I_0_10_add_565_15_lut (.I0(GND_net), .I1(n837[12]), .I2(n699_adj_1363), 
            .I3(n16837), .O(n836_adj_1960[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i455_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n674_adj_1771));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_572_7 (.CI(n16724), .I0(n844_adj_1959[4]), 
            .I1(n328_adj_1894), .CO(n16725));
    SB_LUT4 Q_15__I_0_i488_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n723_adj_1769));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i488_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i33_2_lut (.I0(n19702), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n48));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i33_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY D_15__I_0_10_add_567_13 (.CI(n16805), .I0(n839_adj_1951[10]), 
            .I1(n607_adj_312), .CO(n16806));
    SB_LUT4 add_7655_22_lut (.I0(GND_net), .I1(Product3_mul_temp[22]), .I2(Product4_mul_temp[22]), 
            .I3(n17688), .O(\betaVoltage[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_22 (.CI(n17688), .I0(Product3_mul_temp[22]), .I1(Product4_mul_temp[22]), 
            .CO(n17689));
    SB_LUT4 D_15__I_0_10_add_564_6_lut (.I0(GND_net), .I1(n836_adj_1960[3]), 
            .I2(n255), .I3(n16843), .O(n835_adj_1961[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_566_5 (.CI(n16812), .I0(n838[2]), .I1(n212), 
            .CO(n16813));
    SB_LUT4 add_7655_21_lut (.I0(GND_net), .I1(Product3_mul_temp[21]), .I2(Product4_mul_temp[21]), 
            .I3(n17687), .O(\betaVoltage[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_566_4_lut (.I0(GND_net), .I1(n838[1]), .I2(n163_adj_1898), 
            .I3(n16811), .O(n837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_571_10_lut (.I0(GND_net), .I1(n843[7]), .I2(n478), 
            .I3(n16548), .O(n842[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_572_6_lut (.I0(GND_net), .I1(n844_adj_1959[3]), 
            .I2(n279_adj_314), .I3(n16723), .O(n843_adj_1956[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_6 (.CI(n16723), .I0(n844_adj_1959[3]), 
            .I1(n279_adj_314), .CO(n16724));
    SB_CARRY Q_15__I_0_11_add_568_9 (.CI(n16592), .I0(n840[6]), .I1(n429_c), 
            .CO(n16593));
    SB_LUT4 Q_15__I_0_11_add_568_8_lut (.I0(GND_net), .I1(n840[5]), .I2(n380), 
            .I3(n16591), .O(n839[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_11_lut (.I0(GND_net), .I1(n835[8]), .I2(n527), 
            .I3(n16669), .O(Product2_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_571_9_lut (.I0(GND_net), .I1(n843[6]), .I2(n429_c), 
            .I3(n16547), .O(n842[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_571_8_lut (.I0(GND_net), .I1(n843[5]), .I2(n380), 
            .I3(n16546), .O(n842[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i121_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n178));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i121_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_568_8 (.CI(n16591), .I0(n840[5]), .I1(n380), 
            .CO(n16592));
    SB_LUT4 D_15__I_0_10_add_572_5_lut (.I0(GND_net), .I1(n844_adj_1959[2]), 
            .I2(n230), .I3(n16722), .O(n843_adj_1956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_5 (.CI(n16722), .I0(n844_adj_1959[2]), 
            .I1(n230), .CO(n16723));
    SB_CARRY Q_15__I_0_11_add_571_10 (.CI(n16548), .I0(n843[7]), .I1(n478), 
            .CO(n16549));
    SB_LUT4 D_15__I_0_10_add_572_4_lut (.I0(GND_net), .I1(n844_adj_1959[1]), 
            .I2(n181_adj_1904), .I3(n16721), .O(n843_adj_1956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_570_3_lut (.I0(GND_net), .I1(n842[0]), .I2(n135_c), 
            .I3(n16556), .O(n841_adj_1952[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_4 (.CI(n16721), .I0(n844_adj_1959[1]), 
            .I1(n181_adj_1904), .CO(n16722));
    SB_LUT4 D_15__I_0_10_add_572_3_lut (.I0(GND_net), .I1(n844_adj_1959[0]), 
            .I2(n132_adj_315), .I3(n16720), .O(n843_adj_1956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_568_7_lut (.I0(GND_net), .I1(n840[4]), .I2(n331), 
            .I3(n16590), .O(n839[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_568_7 (.CI(n16590), .I0(n840[4]), .I1(n331), 
            .CO(n16591));
    SB_CARRY Q_15__I_0_11_add_563_11 (.CI(n16669), .I0(n835[8]), .I1(n527), 
            .CO(n16670));
    SB_CARRY Q_15__I_0_11_add_571_8 (.CI(n16546), .I0(n843[5]), .I1(n380), 
            .CO(n16547));
    SB_CARRY D_15__I_0_10_add_572_3 (.CI(n16720), .I0(n844_adj_1959[0]), 
            .I1(n132_adj_315), .CO(n16721));
    SB_CARRY Q_15__I_0_11_add_571_9 (.CI(n16547), .I0(n843[6]), .I1(n429_c), 
            .CO(n16548));
    SB_LUT4 D_15__I_0_10_add_572_2_lut (.I0(GND_net), .I1(n38_adj_316), 
            .I2(n83_adj_317), .I3(GND_net), .O(n843_adj_1956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_572_2 (.CI(GND_net), .I0(n38_adj_316), .I1(n83_adj_317), 
            .CO(n16720));
    SB_CARRY Q_15__I_0_11_add_571_15 (.CI(n16553), .I0(n843[12]), .I1(n723), 
            .CO(n16554));
    SB_LUT4 Q_15__I_0_11_add_563_10_lut (.I0(GND_net), .I1(n835[7]), .I2(n478), 
            .I3(n16668), .O(Product2_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_10 (.CI(n16668), .I0(n835[7]), .I1(n478), 
            .CO(n16669));
    SB_CARRY Q_15__I_0_11_add_564_16 (.CI(n16659), .I0(n836[13]), .I1(n793), 
            .CO(n751_adj_1334));
    SB_LUT4 Q_15__I_0_11_add_563_9_lut (.I0(GND_net), .I1(n835[6]), .I2(n429_c), 
            .I3(n16667), .O(Product2_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_564_14 (.CI(n16657), .I0(n836[11]), .I1(n674), 
            .CO(n16658));
    SB_CARRY Q_15__I_0_11_add_563_9 (.CI(n16667), .I0(n835[6]), .I1(n429_c), 
            .CO(n16668));
    SB_LUT4 Q_15__I_0_11_add_571_15_lut (.I0(GND_net), .I1(n843[12]), .I2(n723), 
            .I3(n16553), .O(n842[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_8_lut (.I0(GND_net), .I1(n835[5]), .I2(n380), 
            .I3(n16666), .O(Product2_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_571_14_lut (.I0(GND_net), .I1(n843[11]), .I2(n674), 
            .I3(n16552), .O(n842[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_8 (.CI(n16666), .I0(n835[5]), .I1(n380), 
            .CO(n16667));
    SB_CARRY Q_15__I_0_11_add_564_15 (.CI(n16658), .I0(n836[12]), .I1(n723), 
            .CO(n16659));
    SB_CARRY Q_15__I_0_11_add_570_3 (.CI(n16556), .I0(n842[0]), .I1(n135_c), 
            .CO(n16557));
    SB_LUT4 D_15__I_0_10_i214_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n316));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i123_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n181));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i123_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i198_2_lut (.I0(\dVoltage[5] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_1317));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i198_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_i247_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n365));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_566_12_lut (.I0(GND_net), .I1(n838_adj_1953[9]), 
            .I2(n576), .I3(n16625), .O(n837_adj_1955[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_12 (.CI(n16625), .I0(n838_adj_1953[9]), 
            .I1(n576), .CO(n16626));
    SB_LUT4 Q_15__I_0_11_add_566_11_lut (.I0(GND_net), .I1(n838_adj_1953[8]), 
            .I2(n527), .I3(n16624), .O(n837_adj_1955[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_11 (.CI(n16624), .I0(n838_adj_1953[8]), 
            .I1(n527), .CO(n16625));
    SB_LUT4 Q_15__I_0_11_add_563_7_lut (.I0(GND_net), .I1(n835[4]), .I2(n331), 
            .I3(n16665), .O(Product2_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i156_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n230_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i222_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n328));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_566_10_lut (.I0(GND_net), .I1(n838_adj_1953[7]), 
            .I2(n478), .I3(n16623), .O(n837_adj_1955[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_i435_2_lut (.I0(\qVoltage[13] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n674));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i435_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i297_2_lut (.I0(\dVoltage[8] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n440_adj_1314));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i297_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY Q_15__I_0_11_add_566_10 (.CI(n16623), .I0(n838_adj_1953[7]), 
            .I1(n478), .CO(n16624));
    SB_LUT4 Q_15__I_0_i255_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n377));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_568_6_lut (.I0(GND_net), .I1(n840[3]), .I2(n282_c), 
            .I3(n16589), .O(n839[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_7 (.CI(n16665), .I0(n835[4]), .I1(n331), 
            .CO(n16666));
    SB_LUT4 Q_15__I_0_i321_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_1757));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i321_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i354_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_1755));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i354_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_299 (.I0(Out_31__N_333), .I1(\preSatVoltage[10] ), 
            .I2(Out_31__N_332), .I3(\Product_mul_temp[26] ), .O(n97));
    defparam i3_4_lut_adj_299.LUT_INIT = 16'h0100;
    SB_CARRY Q_15__I_0_11_add_568_6 (.CI(n16589), .I0(n840[3]), .I1(n282_c), 
            .CO(n16590));
    SB_CARRY D_15__I_0_10_add_566_4 (.CI(n16811), .I0(n838[1]), .I1(n163_adj_1898), 
            .CO(n16812));
    SB_LUT4 Q_15__I_0_11_add_563_6_lut (.I0(GND_net), .I1(n835[3]), .I2(n282_c), 
            .I3(n16664), .O(Product2_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i235_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n347_adj_1751));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_add_573_16_lut (.I0(GND_net), .I1(n845[13]), .I2(n785_adj_318), 
            .I3(n16718), .O(n844_adj_1959[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_16 (.CI(n16718), .I0(n845[13]), .I1(n785_adj_318), 
            .CO(n787_adj_1088));
    SB_LUT4 Q_15__I_0_i453_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n671_adj_1748));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i486_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n720_adj_1746));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i486_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i313_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i313_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Q_15__I_0_11_add_563_6 (.CI(n16664), .I0(n835[3]), .I1(n282_c), 
            .CO(n16665));
    SB_CARRY Q_15__I_0_11_add_564_13 (.CI(n16656), .I0(n836[10]), .I1(n625_c), 
            .CO(n16657));
    SB_LUT4 D_15__I_0_10_add_573_15_lut (.I0(GND_net), .I1(n845[12]), .I2(n723_adj_1912), 
            .I3(n16717), .O(n844_adj_1959[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_11 (.CI(n16549), .I0(n843[8]), .I1(n527), 
            .CO(n16550));
    SB_LUT4 D_15__I_0_i429_2_lut (.I0(\dVoltage[12] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n636_adj_1310));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i429_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY D_15__I_0_10_add_573_15 (.CI(n16717), .I0(n845[12]), .I1(n723_adj_1912), 
            .CO(n16718));
    SB_LUT4 Q_15__I_0_11_add_564_12_lut (.I0(GND_net), .I1(n836[9]), .I2(n576), 
            .I3(n16655), .O(n835[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_i99_2_lut (.I0(\qVoltage[2] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n146));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i99_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_i393_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n582_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i393_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i121_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n178_adj_1736));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i121_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_add_573_14_lut (.I0(GND_net), .I1(n845[11]), .I2(n674_adj_1914), 
            .I3(n16716), .O(n844_adj_1959[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_571_11_lut (.I0(GND_net), .I1(n843[8]), .I2(n527), 
            .I3(n16549), .O(n842[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_21 (.CI(n17687), .I0(Product3_mul_temp[21]), .I1(Product4_mul_temp[21]), 
            .CO(n17688));
    SB_CARRY D_15__I_0_10_add_573_14 (.CI(n16716), .I0(n845[11]), .I1(n674_adj_1914), 
            .CO(n16717));
    SB_LUT4 add_7655_20_lut (.I0(GND_net), .I1(Product3_mul_temp[20]), .I2(Product4_mul_temp[20]), 
            .I3(n17686), .O(\betaVoltage[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_13_lut (.I0(GND_net), .I1(n836[10]), .I2(n625_c), 
            .I3(n16656), .O(n835[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_573_13_lut (.I0(GND_net), .I1(n845[10]), .I2(n625_adj_319), 
            .I3(n16715), .O(n844_adj_1959[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_571_12 (.CI(n16550), .I0(n843[9]), .I1(n576), 
            .CO(n16551));
    SB_CARRY D_15__I_0_10_add_573_13 (.CI(n16715), .I0(n845[10]), .I1(n625_adj_319), 
            .CO(n16716));
    SB_LUT4 Q_15__I_0_11_add_564_14_lut (.I0(GND_net), .I1(n836[11]), .I2(n674), 
            .I3(n16657), .O(n835[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_20 (.CI(n17686), .I0(Product3_mul_temp[20]), .I1(Product4_mul_temp[20]), 
            .CO(n17687));
    SB_LUT4 D_15__I_0_10_add_573_12_lut (.I0(GND_net), .I1(n845[9]), .I2(n576_adj_1918), 
            .I3(n16714), .O(n844_adj_1959[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7655_19_lut (.I0(GND_net), .I1(Product3_mul_temp[19]), .I2(Product4_mul_temp[19]), 
            .I3(n17685), .O(\betaVoltage[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_19 (.CI(n17685), .I0(Product3_mul_temp[19]), .I1(Product4_mul_temp[19]), 
            .CO(n17686));
    SB_LUT4 Q_15__I_0_11_add_571_12_lut (.I0(GND_net), .I1(n843[9]), .I2(n576), 
            .I3(n16550), .O(n842[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_12 (.CI(n16714), .I0(n845[9]), .I1(n576_adj_1918), 
            .CO(n16715));
    SB_CARRY D_15__I_0_10_add_566_13 (.CI(n16820), .I0(n838[10]), .I1(n604_adj_313), 
            .CO(n16821));
    SB_LUT4 Q_15__I_0_11_add_571_16_lut (.I0(GND_net), .I1(n843[13]), .I2(n793), 
            .I3(n16554), .O(n842[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_15_lut (.I0(GND_net), .I1(n836[12]), .I2(n723), 
            .I3(n16658), .O(n835[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_573_11_lut (.I0(GND_net), .I1(n845[8]), .I2(n527_adj_1920), 
            .I3(n16713), .O(n844_adj_1959[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7655_18_lut (.I0(GND_net), .I1(Product3_mul_temp[18]), .I2(Product4_mul_temp[18]), 
            .I3(n17684), .O(\betaVoltage[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_18 (.CI(n17684), .I0(Product3_mul_temp[18]), .I1(Product4_mul_temp[18]), 
            .CO(n17685));
    SB_CARRY Q_15__I_0_11_add_571_13 (.CI(n16551), .I0(n843[10]), .I1(n625_c), 
            .CO(n16552));
    SB_CARRY D_15__I_0_10_add_573_11 (.CI(n16713), .I0(n845[8]), .I1(n527_adj_1920), 
            .CO(n16714));
    SB_LUT4 add_7655_17_lut (.I0(GND_net), .I1(Product3_mul_temp[17]), .I2(Product4_mul_temp[17]), 
            .I3(n17683), .O(\betaVoltage[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_17 (.CI(n17683), .I0(Product3_mul_temp[17]), .I1(Product4_mul_temp[17]), 
            .CO(n17684));
    SB_LUT4 add_7655_16_lut (.I0(GND_net), .I1(Product3_mul_temp[16]), .I2(Product4_mul_temp[16]), 
            .I3(n17682), .O(\Gain1_mul_temp[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_564_16_lut (.I0(GND_net), .I1(n836[13]), .I2(n793), 
            .I3(n16659), .O(n835[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_16 (.CI(n17682), .I0(Product3_mul_temp[16]), .I1(Product4_mul_temp[16]), 
            .CO(n17683));
    SB_LUT4 add_7655_15_lut (.I0(GND_net), .I1(Product3_mul_temp[15]), .I2(Product4_mul_temp[15]), 
            .I3(n17681), .O(\Gain1_mul_temp[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_7655_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7655_15 (.CI(n17681), .I0(Product3_mul_temp[15]), .I1(Product4_mul_temp[15]), 
            .CO(n17682));
    SB_CARRY add_7655_14 (.CI(n17680), .I0(Product3_mul_temp[14]), .I1(Product4_mul_temp[14]), 
            .CO(n17681));
    SB_CARRY add_7655_13 (.CI(n17679), .I0(Product3_mul_temp[13]), .I1(Product4_mul_temp[13]), 
            .CO(n17680));
    SB_CARRY add_7655_12 (.CI(n17678), .I0(Product3_mul_temp[12]), .I1(Product4_mul_temp[12]), 
            .CO(n17679));
    SB_CARRY add_7655_11 (.CI(n17677), .I0(Product3_mul_temp[11]), .I1(Product4_mul_temp[11]), 
            .CO(n17678));
    SB_LUT4 D_15__I_0_10_add_573_10_lut (.I0(GND_net), .I1(n845[7]), .I2(n478_adj_1922), 
            .I3(n16712), .O(n844_adj_1959[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_571_13_lut (.I0(GND_net), .I1(n843[10]), .I2(n625_c), 
            .I3(n16551), .O(n842[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_i346_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i346_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i154_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n227_adj_1734));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i220_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n325_adj_1730));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i220_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n325));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i253_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n374_adj_1728));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i319_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_1724));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i319_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i352_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_1722));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i352_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i253_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n374));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i198_2_lut (.I0(\qVoltage[5] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i198_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY D_15__I_0_10_add_573_10 (.CI(n16712), .I0(n845[7]), .I1(n478_adj_1922), 
            .CO(n16713));
    SB_LUT4 Q_15__I_0_11_i105_2_lut (.I0(\qVoltage[3] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n184));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i72_2_lut (.I0(\qVoltage[2] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n135_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i72_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i138_2_lut (.I0(\qVoltage[4] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n233_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_add_570_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n841_adj_1952[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i451_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n668_adj_1716));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i484_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n717_adj_1714));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i484_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i297_2_lut (.I0(\qVoltage[8] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n440));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i297_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_11_add_563_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(Product2_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_573_9_lut (.I0(GND_net), .I1(n845[6]), .I2(n429_adj_320), 
            .I3(n16711), .O(n844_adj_1959[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_i119_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n175_adj_1704));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i119_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i152_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n224_adj_1702));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_300 (.I0(Out_31__N_332_adj_305), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333_adj_303), .I3(\preSatVoltage[23]_adj_321 ), 
            .O(n19585));
    defparam i1_2_lut_3_lut_4_lut_adj_300.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_11_i336_2_lut (.I0(\qVoltage[10] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i336_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i218_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n322_adj_1698));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i251_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n371_adj_1696));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_301 (.I0(Out_31__N_332_adj_305), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333_adj_303), .I3(\preSatVoltage[19]_adj_322 ), 
            .O(n538_adj_1312));
    defparam i1_2_lut_3_lut_4_lut_adj_301.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_i317_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_1692));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i317_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i350_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_1690));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i350_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_302 (.I0(Out_31__N_332_adj_305), .I1(\Product_mul_temp[26] ), 
            .I2(Out_31__N_333_adj_303), .I3(\preSatVoltage[12]_adj_323 ), 
            .O(n195_adj_1320));
    defparam i1_2_lut_3_lut_4_lut_adj_302.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_11_i429_2_lut (.I0(\qVoltage[12] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n636_adj_1083));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i429_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_i449_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n665_adj_1684));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i482_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n714_adj_1682));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i482_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i319_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i319_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i101_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n148_adj_1673));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i72_2_lut (.I0(\dVoltage[2] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n135_adj_1123));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i72_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i171_2_lut (.I0(\qVoltage[5] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n282_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i204_2_lut (.I0(\qVoltage[6] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n331));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY D_15__I_0_10_add_573_9 (.CI(n16711), .I0(n845[6]), .I1(n429_adj_320), 
            .CO(n16712));
    SB_LUT4 Q_15__I_0_11_add_566_9_lut (.I0(GND_net), .I1(n838_adj_1953[6]), 
            .I2(n429_c), .I3(n16622), .O(n837_adj_1955[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_9 (.CI(n16622), .I0(n838_adj_1953[6]), 
            .I1(n429_c), .CO(n16623));
    SB_LUT4 Q_15__I_0_11_add_566_8_lut (.I0(GND_net), .I1(n838_adj_1953[5]), 
            .I2(n380), .I3(n16621), .O(n837_adj_1955[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_8 (.CI(n16621), .I0(n838_adj_1953[5]), 
            .I1(n380), .CO(n16622));
    SB_LUT4 Q_15__I_0_11_add_566_7_lut (.I0(GND_net), .I1(n838_adj_1953[4]), 
            .I2(n331), .I3(n16620), .O(n837_adj_1955[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_7 (.CI(n16620), .I0(n838_adj_1953[4]), 
            .I1(n331), .CO(n16621));
    SB_LUT4 Q_15__I_0_11_add_566_6_lut (.I0(GND_net), .I1(n838_adj_1953[3]), 
            .I2(n282_c), .I3(n16619), .O(n837_adj_1955[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_6 (.CI(n16619), .I0(n838_adj_1953[3]), 
            .I1(n282_c), .CO(n16620));
    SB_LUT4 Q_15__I_0_11_add_566_5_lut (.I0(GND_net), .I1(n838_adj_1953[2]), 
            .I2(n233_c), .I3(n16618), .O(n837_adj_1955[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_5 (.CI(n16618), .I0(n838_adj_1953[2]), 
            .I1(n233_c), .CO(n16619));
    SB_LUT4 D_15__I_0_10_add_573_8_lut (.I0(GND_net), .I1(n845[5]), .I2(n380_adj_1929), 
            .I3(n16710), .O(n844_adj_1959[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_8 (.CI(n16710), .I0(n845[5]), .I1(n380_adj_1929), 
            .CO(n16711));
    SB_LUT4 D_15__I_0_10_add_573_7_lut (.I0(GND_net), .I1(n845[4]), .I2(n331_adj_1931), 
            .I3(n16709), .O(n844_adj_1959[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_7 (.CI(n16709), .I0(n845[4]), .I1(n331_adj_1931), 
            .CO(n16710));
    SB_LUT4 D_15__I_0_10_add_573_6_lut (.I0(GND_net), .I1(n845[3]), .I2(n282_adj_324), 
            .I3(n16708), .O(n844_adj_1959[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_6 (.CI(n16708), .I0(n845[3]), .I1(n282_adj_324), 
            .CO(n16709));
    SB_LUT4 D_15__I_0_10_add_573_5_lut (.I0(GND_net), .I1(n845[2]), .I2(n233_adj_325), 
            .I3(n16707), .O(n844_adj_1959[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_5 (.CI(n16707), .I0(n845[2]), .I1(n233_adj_325), 
            .CO(n16708));
    SB_LUT4 D_15__I_0_10_add_573_4_lut (.I0(GND_net), .I1(n845[1]), .I2(n184_adj_1935), 
            .I3(n16706), .O(n844_adj_1959[2])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_4 (.CI(n16706), .I0(n845[1]), .I1(n184_adj_1935), 
            .CO(n16707));
    SB_LUT4 Q_15__I_0_11_add_566_4_lut (.I0(GND_net), .I1(n838_adj_1953[1]), 
            .I2(n184), .I3(n16617), .O(n837_adj_1955[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_4 (.CI(n16617), .I0(n838_adj_1953[1]), 
            .I1(n184), .CO(n16618));
    SB_LUT4 Q_15__I_0_11_add_566_3_lut (.I0(GND_net), .I1(n838_adj_1953[0]), 
            .I2(n135_c), .I3(n16616), .O(n837_adj_1955[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_3 (.CI(n16616), .I0(n838_adj_1953[0]), 
            .I1(n135_c), .CO(n16617));
    SB_LUT4 Q_15__I_0_11_add_566_2_lut (.I0(GND_net), .I1(\Product2_mul_temp[2] ), 
            .I2(n86), .I3(GND_net), .O(n837_adj_1955[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_566_2 (.CI(GND_net), .I0(\Product2_mul_temp[2] ), 
            .I1(n86), .CO(n16616));
    SB_LUT4 Q_15__I_0_11_add_567_16_lut (.I0(GND_net), .I1(n839[13]), .I2(n793), 
            .I3(n16614), .O(n838_adj_1953[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_567_16 (.CI(n16614), .I0(n839[13]), .I1(n793), 
            .CO(n763_adj_1331));
    SB_LUT4 Q_15__I_0_11_add_567_15_lut (.I0(GND_net), .I1(n839[12]), .I2(n723), 
            .I3(n16613), .O(n838_adj_1953[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 D_15__I_0_10_add_573_3_lut (.I0(GND_net), .I1(n845[0]), .I2(n135_adj_326), 
            .I3(n16705), .O(n844_adj_1959[1])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_3 (.CI(n16705), .I0(n845[0]), .I1(n135_adj_326), 
            .CO(n16706));
    SB_LUT4 D_15__I_0_10_add_573_2_lut (.I0(GND_net), .I1(n41_adj_327), 
            .I2(n86_adj_328), .I3(GND_net), .O(n844_adj_1959[0])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_573_2 (.CI(GND_net), .I0(n41_adj_327), .I1(n86_adj_328), 
            .CO(n16705));
    SB_LUT4 D_15__I_0_10_add_574_16_lut (.I0(GND_net), .I1(n846[13]), .I2(n789_adj_329), 
            .I3(n16703), .O(n845[14])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_16 (.CI(n16703), .I0(n846[13]), .I1(n789_adj_329), 
            .CO(n791_adj_1086));
    SB_LUT4 D_15__I_0_10_add_574_15_lut (.I0(GND_net), .I1(n846[12]), .I2(n726_adj_1940), 
            .I3(n16702), .O(n845[13])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_15 (.CI(n16702), .I0(n846[12]), .I1(n726_adj_1940), 
            .CO(n16703));
    SB_LUT4 D_15__I_0_10_add_574_14_lut (.I0(GND_net), .I1(n846[11]), .I2(n677_adj_1941), 
            .I3(n16701), .O(n845[12])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_14 (.CI(n16701), .I0(n846[11]), .I1(n677_adj_1941), 
            .CO(n16702));
    SB_LUT4 D_15__I_0_10_i33_2_lut (.I0(n19352), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n48_adj_1670));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i33_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_add_574_13_lut (.I0(GND_net), .I1(n846[10]), .I2(n628_adj_330), 
            .I3(n16700), .O(n845[11])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_13 (.CI(n16700), .I0(n846[10]), .I1(n628_adj_330), 
            .CO(n16701));
    SB_LUT4 D_15__I_0_10_add_574_12_lut (.I0(GND_net), .I1(n846[9]), .I2(n579_adj_1943), 
            .I3(n16699), .O(n845[10])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_12 (.CI(n16699), .I0(n846[9]), .I1(n579_adj_1943), 
            .CO(n16700));
    SB_LUT4 D_15__I_0_10_add_574_11_lut (.I0(GND_net), .I1(n846[8]), .I2(n530_adj_1944), 
            .I3(n16698), .O(n845[9])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_11 (.CI(n16698), .I0(n846[8]), .I1(n530_adj_1944), 
            .CO(n16699));
    SB_LUT4 D_15__I_0_10_add_574_10_lut (.I0(GND_net), .I1(n846[7]), .I2(n481_adj_1945), 
            .I3(n16697), .O(n845[8])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_10 (.CI(n16697), .I0(n846[7]), .I1(n481_adj_1945), 
            .CO(n16698));
    SB_LUT4 D_15__I_0_10_add_574_9_lut (.I0(GND_net), .I1(n846[6]), .I2(n432_adj_331), 
            .I3(n16696), .O(n845[7])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_9 (.CI(n16696), .I0(n846[6]), .I1(n432_adj_331), 
            .CO(n16697));
    SB_LUT4 D_15__I_0_10_add_574_8_lut (.I0(GND_net), .I1(n846[5]), .I2(n383_adj_1947), 
            .I3(n16695), .O(n845[6])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_8 (.CI(n16695), .I0(n846[5]), .I1(n383_adj_1947), 
            .CO(n16696));
    SB_LUT4 D_15__I_0_i105_2_lut (.I0(\dVoltage[3] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n184_adj_1120));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_add_574_7_lut (.I0(GND_net), .I1(n846[4]), .I2(n334_adj_1948), 
            .I3(n16694), .O(n845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_7 (.CI(n16694), .I0(n846[4]), .I1(n334_adj_1948), 
            .CO(n16695));
    SB_LUT4 D_15__I_0_10_add_574_6_lut (.I0(GND_net), .I1(n846[3]), .I2(n285_adj_332), 
            .I3(n16693), .O(n845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY D_15__I_0_10_add_574_6 (.CI(n16693), .I0(n846[3]), .I1(n285_adj_332), 
            .CO(n16694));
    SB_LUT4 D_15__I_0_10_add_574_5_lut (.I0(GND_net), .I1(n846[2]), .I2(n236), 
            .I3(n16692), .O(n845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam D_15__I_0_10_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Q_15__I_0_11_add_563_5_lut (.I0(GND_net), .I1(n835[2]), .I2(n233_c), 
            .I3(n16663), .O(Product2_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_5 (.CI(n16663), .I0(n835[2]), .I1(n233_c), 
            .CO(n16664));
    SB_LUT4 Q_15__I_0_11_add_563_4_lut (.I0(GND_net), .I1(n835[1]), .I2(n184), 
            .I3(n16662), .O(Product2_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Q_15__I_0_11_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Q_15__I_0_11_add_563_4 (.CI(n16662), .I0(n835[1]), .I1(n184), 
            .CO(n16663));
    SB_LUT4 D_15__I_0_i171_2_lut (.I0(\dVoltage[5] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n282_adj_1116));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i301_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_1667));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i301_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i204_2_lut (.I0(\dVoltage[6] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n331_adj_1114));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i237_2_lut (.I0(\dVoltage[7] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n380_adj_1112));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i270_2_lut (.I0(\dVoltage[8] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n429_adj_1110));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i321_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i321_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i371_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n549_adj_1662));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i303_2_lut (.I0(\dVoltage[9] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_1108));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i303_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i210_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n310_adj_1660));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i226_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n334_adj_1948));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i336_2_lut (.I0(\dVoltage[10] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_1106));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i336_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i259_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n383_adj_1947));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i369_2_lut (.I0(\dVoltage[11] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n576_adj_1104));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i402_2_lut (.I0(\dVoltage[12] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n625_adj_1102));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i435_2_lut (.I0(\dVoltage[13] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n674_adj_1101));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i435_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i325_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_1945));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i325_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i468_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n693_adj_1657));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i358_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_1944));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i358_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i468_2_lut (.I0(\dVoltage[14] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n723_adj_1100));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i391_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n579_adj_1943));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i391_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i239_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n353_adj_1655));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i373_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n552_adj_1654));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i457_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n677_adj_1941));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i490_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[13]), 
            .I2(GND_net), .I3(GND_net), .O(n726_adj_1940));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i490_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i208_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n307_adj_1653));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i431_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n638_adj_1649));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i431_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i125_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n184_adj_1935));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i125_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i243_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n359_adj_1648));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i224_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n331_adj_1931));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i443_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n656_adj_1646));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i257_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n380_adj_1929));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i352_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i352_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i385_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n570_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i385_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i117_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n172_adj_1640));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i150_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n221_adj_1638));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i303_2_lut (.I0(\qVoltage[9] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i303_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i451_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n668));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i484_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[10]), 
            .I2(GND_net), .I3(GND_net), .O(n717));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i484_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i3_1_lut (.I0(\Product2_mul_temp[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));
    defparam sub_66_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i4_1_lut (.I0(Product2_mul_temp[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));
    defparam sub_66_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_303 (.I0(Out_31__N_333_adj_303), .I1(\preSatVoltage[10]_adj_304 ), 
            .I2(Out_31__N_332_adj_305), .I3(Look_Up_Table_out1_1[15]), .O(n97_adj_1633));
    defparam i3_4_lut_adj_303.LUT_INIT = 16'h0100;
    SB_LUT4 sub_66_inv_0_i5_1_lut (.I0(Product2_mul_temp[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));
    defparam sub_66_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i6_1_lut (.I0(Product2_mul_temp[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));
    defparam sub_66_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i7_1_lut (.I0(Product2_mul_temp[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));
    defparam sub_66_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i8_1_lut (.I0(Product2_mul_temp[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));
    defparam sub_66_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i9_1_lut (.I0(Product2_mul_temp[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));
    defparam sub_66_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i119_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n175));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i119_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i218_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n322));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i251_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n371));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i10_1_lut (.I0(Product2_mul_temp[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));
    defparam sub_66_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i11_1_lut (.I0(Product2_mul_temp[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));
    defparam sub_66_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i12_1_lut (.I0(Product2_mul_temp[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));
    defparam sub_66_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i13_1_lut (.I0(Product2_mul_temp[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));
    defparam sub_66_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i204_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n301_adj_1629));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i14_1_lut (.I0(Product2_mul_temp[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));
    defparam sub_66_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i317_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i317_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i15_1_lut (.I0(Product2_mul_temp[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));
    defparam sub_66_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i350_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i350_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i237_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[2]), 
            .I2(GND_net), .I3(GND_net), .O(n350_adj_1625));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i383_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n567_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i383_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i449_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n665));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i16_1_lut (.I0(Product2_mul_temp[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));
    defparam sub_66_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i482_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[9]), 
            .I2(GND_net), .I3(GND_net), .O(n714));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i482_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i17_1_lut (.I0(Product2_mul_temp[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));
    defparam sub_66_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i464_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n687_adj_1620));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i18_1_lut (.I0(Product2_mul_temp[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));
    defparam sub_66_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i334_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n494_adj_1618));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i334_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i19_1_lut (.I0(Product2_mul_temp[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));
    defparam sub_66_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i20_1_lut (.I0(Product2_mul_temp[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));
    defparam sub_66_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i437_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n647_adj_1614));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i437_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i21_1_lut (.I0(Product2_mul_temp[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));
    defparam sub_66_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i22_1_lut (.I0(Product2_mul_temp[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));
    defparam sub_66_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i129_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n190));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i129_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i99_2_lut (.I0(\dVoltage[2] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n146_adj_1608));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i99_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 D_15__I_0_10_i241_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[4]), 
            .I2(GND_net), .I3(GND_net), .O(n356_adj_1605));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i23_1_lut (.I0(Product2_mul_temp[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));
    defparam sub_66_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i476_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n705_adj_1600));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i476_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i311_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_1598));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i311_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i24_1_lut (.I0(Product2_mul_temp[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));
    defparam sub_66_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i25_1_lut (.I0(Product2_mul_temp[24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));
    defparam sub_66_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 Q_15__I_0_i216_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n319_adj_1594));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i26_1_lut (.I0(Product2_mul_temp[25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));
    defparam sub_66_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i27_1_lut (.I0(Product2_mul_temp[26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));
    defparam sub_66_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i28_1_lut (.I0(Product2_mul_temp[27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));
    defparam sub_66_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 D_15__I_0_10_i107_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n157_adj_1592));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i117_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n172));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i338_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[3]), 
            .I2(GND_net), .I3(GND_net), .O(n500_adj_1590));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i338_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_66_inv_0_i29_1_lut (.I0(Product2_mul_temp[28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));
    defparam sub_66_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_66_inv_0_i30_1_lut (.I0(Product2_mul_temp[29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));
    defparam sub_66_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 Q_15__I_0_i249_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n368_adj_1577));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i315_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_1573));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i315_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i348_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_1571));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i348_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i216_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n319));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i249_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n368));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i447_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n662_adj_1565));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i480_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n711_adj_1563));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i480_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i309_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_1557));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i309_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i315_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i315_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i323_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_1922));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i323_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i356_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_1920));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i356_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i389_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n576_adj_1918));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i348_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i348_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i115_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n169_adj_1550));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i148_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n218_adj_1546));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i344_2_lut (.I0(\dVoltage[10] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n509_adj_1542));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i344_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i455_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n674_adj_1914));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i214_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n316_adj_1541));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i247_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n365_adj_1539));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i488_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[12]), 
            .I2(GND_net), .I3(GND_net), .O(n723_adj_1912));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i488_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i313_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_1535));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i313_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i381_2_lut (.I0(\dVoltage[11] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n564_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i381_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i346_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_1533));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i346_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i445_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n659_adj_1527));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i478_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n708_adj_1525));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i478_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i478_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n708));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i478_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i123_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n181_adj_1904));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i123_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i111_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n163_adj_1898));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i212_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n313));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i113_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n166_adj_1519));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i447_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n662));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i146_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n215_adj_1517));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i212_2_lut (.I0(\qVoltage[6] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n313_adj_1513));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i480_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[8]), 
            .I2(GND_net), .I3(GND_net), .O(n711));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i480_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i245_2_lut (.I0(\qVoltage[7] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n362));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i459_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n680));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i429_2_lut (.I0(\dVoltage[12] ), .I1(Look_Up_Table_out1_1[15]), 
            .I2(GND_net), .I3(GND_net), .O(n636));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i429_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 Q_15__I_0_i311_2_lut (.I0(\qVoltage[9] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i311_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_304 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[15]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[23] ), .O(n19580));
    defparam i1_2_lut_3_lut_4_lut_adj_304.LUT_INIT = 16'h4044;
    SB_LUT4 Q_15__I_0_i344_2_lut (.I0(\qVoltage[10] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n509));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i344_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i222_2_lut (.I0(\dVoltage[6] ), .I1(Look_Up_Table_out1_1[11]), 
            .I2(GND_net), .I3(GND_net), .O(n328_adj_1894));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i443_2_lut (.I0(\qVoltage[13] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n656));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i476_2_lut (.I0(\qVoltage[14] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n705));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i476_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i245_2_lut (.I0(\dVoltage[7] ), .I1(Look_Up_Table_out1_1[6]), 
            .I2(GND_net), .I3(GND_net), .O(n362_adj_1892));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i441_2_lut (.I0(\dVoltage[13] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n653_adj_1891));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i441_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i299_2_lut (.I0(\dVoltage[9] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_1889));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i299_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i466_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n690_adj_1887));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i466_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i103_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[1]), 
            .I2(GND_net), .I3(GND_net), .O(n151_adj_1886));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_10_i115_2_lut (.I0(\dVoltage[3] ), .I1(Look_Up_Table_out1_1[7]), 
            .I2(GND_net), .I3(GND_net), .O(n169));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_11_i537_2_lut (.I0(\qVoltage[15] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n793));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(61[30:49])
    defparam Q_15__I_0_11_i537_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 D_15__I_0_10_i492_2_lut (.I0(\dVoltage[14] ), .I1(Look_Up_Table_out1_1[14]), 
            .I2(GND_net), .I3(GND_net), .O(n729));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(56[30:49])
    defparam D_15__I_0_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 D_15__I_0_i537_2_lut_2_lut (.I0(\dVoltage[15] ), .I1(\Product_mul_temp[26] ), 
            .I2(GND_net), .I3(GND_net), .O(n793_adj_1098));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(75[30:49])
    defparam D_15__I_0_i537_2_lut_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 Q_15__I_0_i111_2_lut (.I0(\qVoltage[3] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n163));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Q_15__I_0_i144_2_lut (.I0(\qVoltage[4] ), .I1(Look_Up_Table_out1_1[5]), 
            .I2(GND_net), .I3(GND_net), .O(n212_c));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Park_Transform.v(80[30:49])
    defparam Q_15__I_0_i144_2_lut.LUT_INIT = 16'h8888;
    VCC i1 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module Inverse_Clarke_Transform
//

module Inverse_Clarke_Transform (GND_net, \betaVoltage[7] , \betaVoltage[12] , 
            \betaVoltage[3] , \betaVoltage[14] , \betaVoltage[15] , alphaVoltage, 
            \betaVoltage[8] , \betaVoltage[10] , \betaVoltage[5] , \betaVoltage[9] , 
            \betaVoltage[4] , \betaVoltage[13] , \betaVoltage[11] , \Gain1_mul_temp[1] , 
            \Gain1_mul_temp[13] , \Gain1_mul_temp[12] , \Gain1_mul_temp[11] , 
            \Gain1_mul_temp[10] , \Gain1_mul_temp[9] , \Gain1_mul_temp[8] , 
            \Gain1_mul_temp[7] , \Gain1_mul_temp[6] , \Gain1_mul_temp[5] , 
            \Gain1_mul_temp[4] , \Gain1_mul_temp[3] , \betaVoltage[2] , 
            \Gain1_mul_temp[2] , \betaVoltage[6] , \abcVoltage_1[31] , 
            \abcVoltage_1[30] , \abcVoltage_1[29] , \abcVoltage_1[28] , 
            \abcVoltage_1[27] , \abcVoltage_1[26] , \abcVoltage_1[25] , 
            \abcVoltage_1[24] , \abcVoltage_1[23] , \abcVoltage_1[22] , 
            \abcVoltage_1[21] , \abcVoltage_1[20] , \abcVoltage_1[19] , 
            \abcVoltage_1[18] , \abcVoltage_1[17] , \abcVoltage_1[16] , 
            \abcVoltage_1[15] , \abcVoltage_1[14] , \abcVoltage_2[31] , 
            \abcVoltage_2[30] , \abcVoltage_2[29] , \abcVoltage_2[28] , 
            \abcVoltage_2[27] , \abcVoltage_2[26] , \abcVoltage_2[25] , 
            \abcVoltage_2[24] , \abcVoltage_2[23] , \abcVoltage_2[22] , 
            \abcVoltage_2[21] , \abcVoltage_2[20] , \abcVoltage_2[19] , 
            \abcVoltage_2[18] , \abcVoltage_2[17] , \abcVoltage_2[16] , 
            \abcVoltage_2[15] , \abcVoltage_2[14] , \abcVoltage_2[13] , 
            \abcVoltage_2[12] , \abcVoltage_2[11] , \abcVoltage_2[10] , 
            \abcVoltage_2[9] , \abcVoltage_2[8] , \abcVoltage_2[7] , \abcVoltage_2[6] , 
            \abcVoltage_2[5] , \abcVoltage_2[4] , \abcVoltage_2[3] , \abcVoltage_2[2] , 
            \abcVoltage_2[1] ) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \betaVoltage[7] ;
    input \betaVoltage[12] ;
    input \betaVoltage[3] ;
    input \betaVoltage[14] ;
    input \betaVoltage[15] ;
    input [15:0]alphaVoltage;
    input \betaVoltage[8] ;
    input \betaVoltage[10] ;
    input \betaVoltage[5] ;
    input \betaVoltage[9] ;
    input \betaVoltage[4] ;
    input \betaVoltage[13] ;
    input \betaVoltage[11] ;
    input \Gain1_mul_temp[1] ;
    output \Gain1_mul_temp[13] ;
    output \Gain1_mul_temp[12] ;
    output \Gain1_mul_temp[11] ;
    output \Gain1_mul_temp[10] ;
    output \Gain1_mul_temp[9] ;
    output \Gain1_mul_temp[8] ;
    output \Gain1_mul_temp[7] ;
    output \Gain1_mul_temp[6] ;
    output \Gain1_mul_temp[5] ;
    output \Gain1_mul_temp[4] ;
    output \Gain1_mul_temp[3] ;
    input \betaVoltage[2] ;
    input \Gain1_mul_temp[2] ;
    input \betaVoltage[6] ;
    output \abcVoltage_1[31] ;
    output \abcVoltage_1[30] ;
    output \abcVoltage_1[29] ;
    output \abcVoltage_1[28] ;
    output \abcVoltage_1[27] ;
    output \abcVoltage_1[26] ;
    output \abcVoltage_1[25] ;
    output \abcVoltage_1[24] ;
    output \abcVoltage_1[23] ;
    output \abcVoltage_1[22] ;
    output \abcVoltage_1[21] ;
    output \abcVoltage_1[20] ;
    output \abcVoltage_1[19] ;
    output \abcVoltage_1[18] ;
    output \abcVoltage_1[17] ;
    output \abcVoltage_1[16] ;
    output \abcVoltage_1[15] ;
    output \abcVoltage_1[14] ;
    output \abcVoltage_2[31] ;
    output \abcVoltage_2[30] ;
    output \abcVoltage_2[29] ;
    output \abcVoltage_2[28] ;
    output \abcVoltage_2[27] ;
    output \abcVoltage_2[26] ;
    output \abcVoltage_2[25] ;
    output \abcVoltage_2[24] ;
    output \abcVoltage_2[23] ;
    output \abcVoltage_2[22] ;
    output \abcVoltage_2[21] ;
    output \abcVoltage_2[20] ;
    output \abcVoltage_2[19] ;
    output \abcVoltage_2[18] ;
    output \abcVoltage_2[17] ;
    output \abcVoltage_2[16] ;
    output \abcVoltage_2[15] ;
    output \abcVoltage_2[14] ;
    output \abcVoltage_2[13] ;
    output \abcVoltage_2[12] ;
    output \abcVoltage_2[11] ;
    output \abcVoltage_2[10] ;
    output \abcVoltage_2[9] ;
    output \abcVoltage_2[8] ;
    output \abcVoltage_2[7] ;
    output \abcVoltage_2[6] ;
    output \abcVoltage_2[5] ;
    output \abcVoltage_2[4] ;
    output \abcVoltage_2[3] ;
    output \abcVoltage_2[2] ;
    output \abcVoltage_2[1] ;
    
    wire [14:0]n839;
    wire [14:0]n840;
    
    wire n15602, n15603, n15601, n15600, n15599;
    wire [14:0]n844;
    wire [14:0]n845;
    
    wire n15481, n15832;
    wire [14:0]n836;
    
    wire n15833;
    wire [13:0]n7479;
    
    wire n17703;
    wire [14:0]n835;
    
    wire n15831, n17704, n15482, n15480, n17702, n17701, n15479;
    wire [17:0]n1;
    
    wire n17700, n17699, n17698, n17697, n15598, n15478, n15477, 
        n15476, n15475, n15474, n15473, n15472;
    wire [14:0]n841;
    
    wire n15566, n771, n15565, n15564, n15563, n15562, n15561, 
        n15560, n15559, n15558, n15557, n15556, n15555, n15606, 
        n15607, n15605;
    wire [14:0]n842;
    
    wire n15522, n15834, n775, n15521, n15520, n15519;
    wire [14:0]n837;
    
    wire n15829, n15518, n15517, n755, n15516, n15828, n15515, 
        n15514;
    wire [33:0]Add1_cast_1;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Clarke_Transform.v(46[22:33])
    
    wire n15972, n15971, n15970, n15513, n15969, n15968, n15604, 
        n15967, n15512, n18410, n791, n18409, n18408, n18407, 
        n18406, n18405, n18404, n18403, n18402, n18401, n18400, 
        n18399;
    wire [31:0]Gain1_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Clarke_Transform.v(37[22:36])
    
    wire n18398, n7494, n18397, n787, n18396, n783, n18395;
    wire [14:0]n843;
    
    wire n779, n18394, n18393, n18392, n767, n18391, n763, n18390;
    wire [14:0]n838;
    
    wire n759, n18389, n18388, n751, n18387, n747, n18386;
    wire [14:0]n834;
    
    wire n743, n18385;
    wire [14:0]n833;
    
    wire n739, n18384;
    wire [14:0]n832;
    
    wire n15966, n15965, n15511, n17709, n17708, n17707, n15964, 
        n15963, n15509, n15962, n15961, n15827, n15960, n15508, 
        n15959, n15507;
    wire [33:0]n1_adj_1007;
    
    wire n15958, n15957, VCC_net, n15506, n15505, n15504, n15503, 
        n15502, n15501, n15500, n15499, n15498, n15496, n15495, 
        n15494, n15493, n15492, n15491, n15490, n15489, n15488, 
        n15826, n15487, n15486, n15485, n15483, n15881, n15880, 
        n15879, n15878, n15877, n15876, n15875, n15874, n15873, 
        n15872, n15871, n15870, n15868, n15867, n15866, n15865, 
        n15864, n15863, n15862, n15861, n15860, n15859, n15858, 
        n15857, n15855, n15854, n15853, n15852, n15851, n15850, 
        n15849, n15848, n15847, n15846, n15845, n15844, n15842, 
        n15841, n15840, n15839, n15838, n15825, n15824, n15823, 
        n15822, n15821, n15820, n17706, n17705, n15819, n15818, 
        n15816, n15815, n15814, n15813, n15812, n15811, n15810, 
        n15809, n15808, n15807, n15837, n15806, n15805, n15836, 
        n15835, n15719, n15718, n15717, n15716, n15608, n15715, 
        n15714, n15713, n15712, n15711, n15710, n15709, n15708, 
        n15707, n15622, n15706, n15705, n15621, n15704, n15703;
    wire [31:0]n1_adj_1008;
    
    wire n15702, n15701, n15700, n15699, n15698, n15697, n15696, 
        n15695, n15694, n15693, n15692, n15691, n15690, n15689, 
        n15688, n15687, n15686, n15685, n15684, n15683, n15682, 
        n15681, n15680, n15679, n15678, n15620, n15619, n15618, 
        n15617, n15616, n15677, n15615, n15676, n15675, n15614, 
        n15674, n15673, n15613, n15672, n15612, n15611, n15609;
    
    SB_LUT4 Beta_15__I_0_add_568_7_lut (.I0(GND_net), .I1(n840[6]), .I2(GND_net), 
            .I3(n15602), .O(n839[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_7 (.CI(n15602), .I0(n840[6]), .I1(GND_net), 
            .CO(n15603));
    SB_LUT4 Beta_15__I_0_add_568_6_lut (.I0(GND_net), .I1(n840[5]), .I2(\betaVoltage[7] ), 
            .I3(n15601), .O(n839[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_6 (.CI(n15601), .I0(n840[5]), .I1(\betaVoltage[7] ), 
            .CO(n15602));
    SB_LUT4 Beta_15__I_0_add_568_5_lut (.I0(GND_net), .I1(n840[4]), .I2(\betaVoltage[7] ), 
            .I3(n15600), .O(n839[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_5 (.CI(n15600), .I0(n840[4]), .I1(\betaVoltage[7] ), 
            .CO(n15601));
    SB_LUT4 Beta_15__I_0_add_568_4_lut (.I0(GND_net), .I1(n840[3]), .I2(GND_net), 
            .I3(n15599), .O(n839[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_573_12_lut (.I0(GND_net), .I1(n845[11]), .I2(\betaVoltage[12] ), 
            .I3(n15481), .O(n844[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_4 (.CI(n15832), .I0(n836[3]), .I1(GND_net), 
            .CO(n15833));
    SB_LUT4 add_5933_9_lut (.I0(GND_net), .I1(GND_net), .I2(GND_net), 
            .I3(n17703), .O(n7479[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_4 (.CI(n15599), .I0(n840[3]), .I1(GND_net), 
            .CO(n15600));
    SB_LUT4 Beta_15__I_0_add_564_3_lut (.I0(GND_net), .I1(n836[2]), .I2(\betaVoltage[3] ), 
            .I3(n15831), .O(n835[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_9 (.CI(n17703), .I0(GND_net), .I1(GND_net), .CO(n17704));
    SB_CARRY Beta_15__I_0_add_573_12 (.CI(n15481), .I0(n845[11]), .I1(\betaVoltage[12] ), 
            .CO(n15482));
    SB_LUT4 Beta_15__I_0_add_573_11_lut (.I0(GND_net), .I1(n845[10]), .I2(GND_net), 
            .I3(n15480), .O(n844[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5933_8_lut (.I0(GND_net), .I1(GND_net), .I2(\betaVoltage[14] ), 
            .I3(n17702), .O(n7479[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_11 (.CI(n15480), .I0(n845[10]), .I1(GND_net), 
            .CO(n15481));
    SB_CARRY add_5933_8 (.CI(n17702), .I0(GND_net), .I1(\betaVoltage[14] ), 
            .CO(n17703));
    SB_LUT4 add_5933_7_lut (.I0(GND_net), .I1(\betaVoltage[15] ), .I2(\betaVoltage[14] ), 
            .I3(n17701), .O(n7479[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_573_10_lut (.I0(GND_net), .I1(n845[9]), .I2(\betaVoltage[12] ), 
            .I3(n15479), .O(n844[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_10 (.CI(n15479), .I0(n845[9]), .I1(\betaVoltage[12] ), 
            .CO(n15480));
    SB_CARRY add_5933_7 (.CI(n17701), .I0(\betaVoltage[15] ), .I1(\betaVoltage[14] ), 
            .CO(n17702));
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(alphaVoltage[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5933_6_lut (.I0(GND_net), .I1(GND_net), .I2(GND_net), 
            .I3(n17700), .O(n7479[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_6 (.CI(n17700), .I0(GND_net), .I1(GND_net), .CO(n17701));
    SB_LUT4 add_5933_5_lut (.I0(GND_net), .I1(GND_net), .I2(\betaVoltage[14] ), 
            .I3(n17699), .O(n7479[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_5 (.CI(n17699), .I0(GND_net), .I1(\betaVoltage[14] ), 
            .CO(n17700));
    SB_LUT4 add_5933_4_lut (.I0(GND_net), .I1(\betaVoltage[15] ), .I2(\betaVoltage[14] ), 
            .I3(n17698), .O(n7479[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_4 (.CI(n17698), .I0(\betaVoltage[15] ), .I1(\betaVoltage[14] ), 
            .CO(n17699));
    SB_LUT4 add_5933_3_lut (.I0(GND_net), .I1(GND_net), .I2(GND_net), 
            .I3(n17697), .O(n7479[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_3 (.CI(n17697), .I0(GND_net), .I1(GND_net), .CO(n17698));
    SB_LUT4 Beta_15__I_0_add_568_3_lut (.I0(GND_net), .I1(n840[2]), .I2(\betaVoltage[7] ), 
            .I3(n15598), .O(n839[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5933_2_lut (.I0(GND_net), .I1(\betaVoltage[15] ), .I2(\betaVoltage[14] ), 
            .I3(GND_net), .O(n7479[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_2 (.CI(GND_net), .I0(\betaVoltage[15] ), .I1(\betaVoltage[14] ), 
            .CO(n17697));
    SB_LUT4 Beta_15__I_0_add_573_9_lut (.I0(GND_net), .I1(n845[8]), .I2(\betaVoltage[12] ), 
            .I3(n15478), .O(n844[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_9 (.CI(n15478), .I0(n845[8]), .I1(\betaVoltage[12] ), 
            .CO(n15479));
    SB_LUT4 Beta_15__I_0_add_573_8_lut (.I0(GND_net), .I1(n845[7]), .I2(\betaVoltage[12] ), 
            .I3(n15477), .O(n844[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_8 (.CI(n15477), .I0(n845[7]), .I1(\betaVoltage[12] ), 
            .CO(n15478));
    SB_LUT4 Beta_15__I_0_add_573_7_lut (.I0(GND_net), .I1(n845[6]), .I2(GND_net), 
            .I3(n15476), .O(n844[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_7 (.CI(n15476), .I0(n845[6]), .I1(GND_net), 
            .CO(n15477));
    SB_LUT4 Beta_15__I_0_add_573_6_lut (.I0(GND_net), .I1(n845[5]), .I2(\betaVoltage[12] ), 
            .I3(n15475), .O(n844[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_6 (.CI(n15475), .I0(n845[5]), .I1(\betaVoltage[12] ), 
            .CO(n15476));
    SB_LUT4 Beta_15__I_0_add_573_5_lut (.I0(GND_net), .I1(n845[4]), .I2(\betaVoltage[12] ), 
            .I3(n15474), .O(n844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_5 (.CI(n15474), .I0(n845[4]), .I1(\betaVoltage[12] ), 
            .CO(n15475));
    SB_LUT4 Beta_15__I_0_add_573_4_lut (.I0(GND_net), .I1(n845[3]), .I2(GND_net), 
            .I3(n15473), .O(n844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_4 (.CI(n15473), .I0(n845[3]), .I1(GND_net), 
            .CO(n15474));
    SB_LUT4 Beta_15__I_0_add_573_3_lut (.I0(GND_net), .I1(n845[2]), .I2(\betaVoltage[12] ), 
            .I3(n15472), .O(n844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_3 (.CI(n15472), .I0(n845[2]), .I1(\betaVoltage[12] ), 
            .CO(n15473));
    SB_LUT4 Beta_15__I_0_add_573_2_lut (.I0(GND_net), .I1(n7479[0]), .I2(\betaVoltage[12] ), 
            .I3(GND_net), .O(n844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_569_14_lut (.I0(GND_net), .I1(n841[13]), .I2(GND_net), 
            .I3(n15566), .O(n840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_14 (.CI(n15566), .I0(n841[13]), .I1(GND_net), 
            .CO(n771));
    SB_LUT4 Beta_15__I_0_add_569_13_lut (.I0(GND_net), .I1(n841[12]), .I2(\betaVoltage[8] ), 
            .I3(n15565), .O(n840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_13 (.CI(n15565), .I0(n841[12]), .I1(\betaVoltage[8] ), 
            .CO(n15566));
    SB_LUT4 Beta_15__I_0_add_569_12_lut (.I0(GND_net), .I1(n841[11]), .I2(\betaVoltage[8] ), 
            .I3(n15564), .O(n840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_12 (.CI(n15564), .I0(n841[11]), .I1(\betaVoltage[8] ), 
            .CO(n15565));
    SB_LUT4 Beta_15__I_0_add_569_11_lut (.I0(GND_net), .I1(n841[10]), .I2(GND_net), 
            .I3(n15563), .O(n840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_11 (.CI(n15563), .I0(n841[10]), .I1(GND_net), 
            .CO(n15564));
    SB_LUT4 Beta_15__I_0_add_569_10_lut (.I0(GND_net), .I1(n841[9]), .I2(\betaVoltage[8] ), 
            .I3(n15562), .O(n840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_10 (.CI(n15562), .I0(n841[9]), .I1(\betaVoltage[8] ), 
            .CO(n15563));
    SB_LUT4 Beta_15__I_0_add_569_9_lut (.I0(GND_net), .I1(n841[8]), .I2(\betaVoltage[8] ), 
            .I3(n15561), .O(n840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_9 (.CI(n15561), .I0(n841[8]), .I1(\betaVoltage[8] ), 
            .CO(n15562));
    SB_LUT4 Beta_15__I_0_add_569_8_lut (.I0(GND_net), .I1(n841[7]), .I2(\betaVoltage[8] ), 
            .I3(n15560), .O(n840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_8 (.CI(n15560), .I0(n841[7]), .I1(\betaVoltage[8] ), 
            .CO(n15561));
    SB_LUT4 Beta_15__I_0_add_569_7_lut (.I0(GND_net), .I1(n841[6]), .I2(GND_net), 
            .I3(n15559), .O(n840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_7 (.CI(n15559), .I0(n841[6]), .I1(GND_net), 
            .CO(n15560));
    SB_LUT4 Beta_15__I_0_add_569_6_lut (.I0(GND_net), .I1(n841[5]), .I2(\betaVoltage[8] ), 
            .I3(n15558), .O(n840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_6 (.CI(n15558), .I0(n841[5]), .I1(\betaVoltage[8] ), 
            .CO(n15559));
    SB_LUT4 Beta_15__I_0_add_569_5_lut (.I0(GND_net), .I1(n841[4]), .I2(\betaVoltage[8] ), 
            .I3(n15557), .O(n840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_5 (.CI(n15557), .I0(n841[4]), .I1(\betaVoltage[8] ), 
            .CO(n15558));
    SB_LUT4 Beta_15__I_0_add_569_4_lut (.I0(GND_net), .I1(n841[3]), .I2(GND_net), 
            .I3(n15556), .O(n840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_4 (.CI(n15556), .I0(n841[3]), .I1(GND_net), 
            .CO(n15557));
    SB_LUT4 Beta_15__I_0_add_569_3_lut (.I0(GND_net), .I1(n841[2]), .I2(\betaVoltage[8] ), 
            .I3(n15555), .O(n840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_3 (.CI(n15555), .I0(n841[2]), .I1(\betaVoltage[8] ), 
            .CO(n15556));
    SB_LUT4 Beta_15__I_0_add_569_2_lut (.I0(GND_net), .I1(\betaVoltage[10] ), 
            .I2(\betaVoltage[8] ), .I3(GND_net), .O(n840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_569_2 (.CI(GND_net), .I0(\betaVoltage[10] ), 
            .I1(\betaVoltage[8] ), .CO(n15555));
    SB_CARRY Beta_15__I_0_add_568_11 (.CI(n15606), .I0(n840[10]), .I1(GND_net), 
            .CO(n15607));
    SB_CARRY Beta_15__I_0_add_564_3 (.CI(n15831), .I0(n836[2]), .I1(\betaVoltage[3] ), 
            .CO(n15832));
    SB_LUT4 Beta_15__I_0_add_568_10_lut (.I0(GND_net), .I1(n840[9]), .I2(\betaVoltage[7] ), 
            .I3(n15605), .O(n839[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_2_lut (.I0(GND_net), .I1(\betaVoltage[5] ), 
            .I2(\betaVoltage[3] ), .I3(GND_net), .O(n835[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_3 (.CI(n15598), .I0(n840[2]), .I1(\betaVoltage[7] ), 
            .CO(n15599));
    SB_LUT4 Beta_15__I_0_add_568_2_lut (.I0(GND_net), .I1(\betaVoltage[9] ), 
            .I2(\betaVoltage[7] ), .I3(GND_net), .O(n839[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_570_14_lut (.I0(GND_net), .I1(n842[13]), .I2(GND_net), 
            .I3(n15522), .O(n841[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_2 (.CI(GND_net), .I0(\betaVoltage[9] ), 
            .I1(\betaVoltage[7] ), .CO(n15598));
    SB_CARRY Beta_15__I_0_add_564_5 (.CI(n15833), .I0(n836[4]), .I1(\betaVoltage[3] ), 
            .CO(n15834));
    SB_CARRY Beta_15__I_0_add_570_14 (.CI(n15522), .I0(n842[13]), .I1(GND_net), 
            .CO(n775));
    SB_LUT4 Beta_15__I_0_add_570_13_lut (.I0(GND_net), .I1(n842[12]), .I2(\betaVoltage[9] ), 
            .I3(n15521), .O(n841[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_13 (.CI(n15521), .I0(n842[12]), .I1(\betaVoltage[9] ), 
            .CO(n15522));
    SB_LUT4 Beta_15__I_0_add_570_12_lut (.I0(GND_net), .I1(n842[11]), .I2(\betaVoltage[9] ), 
            .I3(n15520), .O(n841[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_12 (.CI(n15520), .I0(n842[11]), .I1(\betaVoltage[9] ), 
            .CO(n15521));
    SB_LUT4 Beta_15__I_0_add_570_11_lut (.I0(GND_net), .I1(n842[10]), .I2(GND_net), 
            .I3(n15519), .O(n841[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_2 (.CI(GND_net), .I0(\betaVoltage[5] ), 
            .I1(\betaVoltage[3] ), .CO(n15831));
    SB_LUT4 Beta_15__I_0_add_565_14_lut (.I0(GND_net), .I1(n837[13]), .I2(GND_net), 
            .I3(n15829), .O(n836[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_11 (.CI(n15519), .I0(n842[10]), .I1(GND_net), 
            .CO(n15520));
    SB_LUT4 Beta_15__I_0_add_570_10_lut (.I0(GND_net), .I1(n842[9]), .I2(\betaVoltage[9] ), 
            .I3(n15518), .O(n841[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_10 (.CI(n15518), .I0(n842[9]), .I1(\betaVoltage[9] ), 
            .CO(n15519));
    SB_LUT4 Beta_15__I_0_add_570_9_lut (.I0(GND_net), .I1(n842[8]), .I2(\betaVoltage[9] ), 
            .I3(n15517), .O(n841[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_14 (.CI(n15829), .I0(n837[13]), .I1(GND_net), 
            .CO(n755));
    SB_CARRY Beta_15__I_0_add_570_9 (.CI(n15517), .I0(n842[8]), .I1(\betaVoltage[9] ), 
            .CO(n15518));
    SB_LUT4 Beta_15__I_0_add_570_8_lut (.I0(GND_net), .I1(n842[7]), .I2(\betaVoltage[9] ), 
            .I3(n15516), .O(n841[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_565_13_lut (.I0(GND_net), .I1(n837[12]), .I2(\betaVoltage[4] ), 
            .I3(n15828), .O(n836[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_8 (.CI(n15516), .I0(n842[7]), .I1(\betaVoltage[9] ), 
            .CO(n15517));
    SB_LUT4 Beta_15__I_0_add_570_7_lut (.I0(GND_net), .I1(n842[6]), .I2(GND_net), 
            .I3(n15515), .O(n841[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_7 (.CI(n15515), .I0(n842[6]), .I1(GND_net), 
            .CO(n15516));
    SB_LUT4 sub_67_inv_0_i12_1_lut (.I0(alphaVoltage[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));
    defparam sub_67_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i13_1_lut (.I0(alphaVoltage[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));
    defparam sub_67_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i14_1_lut (.I0(alphaVoltage[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));
    defparam sub_67_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i15_1_lut (.I0(alphaVoltage[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));
    defparam sub_67_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i16_1_lut (.I0(alphaVoltage[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));
    defparam sub_67_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 Beta_15__I_0_add_570_6_lut (.I0(GND_net), .I1(n842[5]), .I2(\betaVoltage[9] ), 
            .I3(n15514), .O(n841[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n15972), .O(Add1_cast_1[32])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n15971), .O(Add1_cast_1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_17 (.CI(n15971), .I0(GND_net), .I1(n1[15]), 
            .CO(n15972));
    SB_CARRY Beta_15__I_0_add_568_10 (.CI(n15605), .I0(n840[9]), .I1(\betaVoltage[7] ), 
            .CO(n15606));
    SB_CARRY Beta_15__I_0_add_565_13 (.CI(n15828), .I0(n837[12]), .I1(\betaVoltage[4] ), 
            .CO(n15829));
    SB_LUT4 Alpha_15__I_0_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n15970), .O(Add1_cast_1[30])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_6 (.CI(n15514), .I0(n842[5]), .I1(\betaVoltage[9] ), 
            .CO(n15515));
    SB_CARRY Alpha_15__I_0_add_3_16 (.CI(n15970), .I0(GND_net), .I1(n1[14]), 
            .CO(n15971));
    SB_LUT4 Beta_15__I_0_add_570_5_lut (.I0(GND_net), .I1(n842[4]), .I2(\betaVoltage[9] ), 
            .I3(n15513), .O(n841[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n15969), .O(Add1_cast_1[29])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_15 (.CI(n15969), .I0(GND_net), .I1(n1[13]), 
            .CO(n15970));
    SB_LUT4 Alpha_15__I_0_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n15968), .O(Add1_cast_1[28])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_9_lut (.I0(GND_net), .I1(n840[8]), .I2(\betaVoltage[7] ), 
            .I3(n15604), .O(n839[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_14 (.CI(n15968), .I0(GND_net), .I1(n1[12]), 
            .CO(n15969));
    SB_LUT4 Alpha_15__I_0_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n15967), .O(Add1_cast_1[27])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_5 (.CI(n15513), .I0(n842[4]), .I1(\betaVoltage[9] ), 
            .CO(n15514));
    SB_LUT4 Beta_15__I_0_add_570_4_lut (.I0(GND_net), .I1(n842[3]), .I2(GND_net), 
            .I3(n15512), .O(n841[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_4 (.CI(n15512), .I0(n842[3]), .I1(GND_net), 
            .CO(n15513));
    SB_CARRY Alpha_15__I_0_add_3_13 (.CI(n15967), .I0(GND_net), .I1(n1[11]), 
            .CO(n15968));
    SB_LUT4 Beta_15__I_0_add_574_14_lut (.I0(GND_net), .I1(n7479[13]), .I2(GND_net), 
            .I3(n18410), .O(n845[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_14 (.CI(n18410), .I0(n7479[13]), .I1(GND_net), 
            .CO(n791));
    SB_LUT4 Beta_15__I_0_add_574_13_lut (.I0(GND_net), .I1(n7479[12]), .I2(\betaVoltage[13] ), 
            .I3(n18409), .O(n845[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_13 (.CI(n18409), .I0(n7479[12]), .I1(\betaVoltage[13] ), 
            .CO(n18410));
    SB_LUT4 Beta_15__I_0_add_574_12_lut (.I0(GND_net), .I1(n7479[11]), .I2(\betaVoltage[13] ), 
            .I3(n18408), .O(n845[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_12 (.CI(n18408), .I0(n7479[11]), .I1(\betaVoltage[13] ), 
            .CO(n18409));
    SB_LUT4 Beta_15__I_0_add_574_11_lut (.I0(GND_net), .I1(n7479[10]), .I2(GND_net), 
            .I3(n18407), .O(n845[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_11 (.CI(n18407), .I0(n7479[10]), .I1(GND_net), 
            .CO(n18408));
    SB_LUT4 Beta_15__I_0_add_574_10_lut (.I0(GND_net), .I1(n7479[9]), .I2(\betaVoltage[13] ), 
            .I3(n18406), .O(n845[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_10 (.CI(n18406), .I0(n7479[9]), .I1(\betaVoltage[13] ), 
            .CO(n18407));
    SB_LUT4 Beta_15__I_0_add_574_9_lut (.I0(GND_net), .I1(n7479[8]), .I2(\betaVoltage[13] ), 
            .I3(n18405), .O(n845[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_9 (.CI(n18405), .I0(n7479[8]), .I1(\betaVoltage[13] ), 
            .CO(n18406));
    SB_LUT4 Beta_15__I_0_add_574_8_lut (.I0(GND_net), .I1(n7479[7]), .I2(\betaVoltage[13] ), 
            .I3(n18404), .O(n845[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_8 (.CI(n18404), .I0(n7479[7]), .I1(\betaVoltage[13] ), 
            .CO(n18405));
    SB_LUT4 Beta_15__I_0_add_574_7_lut (.I0(GND_net), .I1(n7479[6]), .I2(GND_net), 
            .I3(n18403), .O(n845[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_7 (.CI(n18403), .I0(n7479[6]), .I1(GND_net), 
            .CO(n18404));
    SB_LUT4 Beta_15__I_0_add_574_6_lut (.I0(GND_net), .I1(n7479[5]), .I2(\betaVoltage[13] ), 
            .I3(n18402), .O(n845[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_6 (.CI(n18402), .I0(n7479[5]), .I1(\betaVoltage[13] ), 
            .CO(n18403));
    SB_LUT4 Beta_15__I_0_add_574_5_lut (.I0(GND_net), .I1(n7479[4]), .I2(\betaVoltage[13] ), 
            .I3(n18401), .O(n845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_5 (.CI(n18401), .I0(n7479[4]), .I1(\betaVoltage[13] ), 
            .CO(n18402));
    SB_LUT4 Beta_15__I_0_add_574_4_lut (.I0(GND_net), .I1(n7479[3]), .I2(GND_net), 
            .I3(n18400), .O(n845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_4 (.CI(n18400), .I0(n7479[3]), .I1(GND_net), 
            .CO(n18401));
    SB_LUT4 Beta_15__I_0_add_574_3_lut (.I0(GND_net), .I1(n7479[2]), .I2(\betaVoltage[13] ), 
            .I3(n18399), .O(n845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_3 (.CI(n18399), .I0(n7479[2]), .I1(\betaVoltage[13] ), 
            .CO(n18400));
    SB_LUT4 Beta_15__I_0_add_574_2_lut (.I0(GND_net), .I1(n7479[1]), .I2(\betaVoltage[13] ), 
            .I3(GND_net), .O(n845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_574_2 (.CI(GND_net), .I0(n7479[1]), .I1(\betaVoltage[13] ), 
            .CO(n18399));
    SB_LUT4 add_1225_17_lut (.I0(GND_net), .I1(\betaVoltage[15] ), .I2(GND_net), 
            .I3(n18398), .O(Gain1_mul_temp[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1225_16_lut (.I0(GND_net), .I1(n7494), .I2(n791), .I3(n18397), 
            .O(Gain1_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_16 (.CI(n18397), .I0(n7494), .I1(n791), .CO(n18398));
    SB_LUT4 add_1225_15_lut (.I0(GND_net), .I1(n845[14]), .I2(n787), .I3(n18396), 
            .O(Gain1_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_15 (.CI(n18396), .I0(n845[14]), .I1(n787), .CO(n18397));
    SB_LUT4 add_1225_14_lut (.I0(GND_net), .I1(n844[14]), .I2(n783), .I3(n18395), 
            .O(Gain1_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_14 (.CI(n18395), .I0(n844[14]), .I1(n783), .CO(n18396));
    SB_LUT4 add_1225_13_lut (.I0(GND_net), .I1(n843[14]), .I2(n779), .I3(n18394), 
            .O(Gain1_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_13 (.CI(n18394), .I0(n843[14]), .I1(n779), .CO(n18395));
    SB_LUT4 add_1225_12_lut (.I0(GND_net), .I1(n842[14]), .I2(n775), .I3(n18393), 
            .O(Gain1_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_12 (.CI(n18393), .I0(n842[14]), .I1(n775), .CO(n18394));
    SB_LUT4 add_1225_11_lut (.I0(GND_net), .I1(n841[14]), .I2(n771), .I3(n18392), 
            .O(Gain1_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_11 (.CI(n18392), .I0(n841[14]), .I1(n771), .CO(n18393));
    SB_LUT4 add_1225_10_lut (.I0(GND_net), .I1(n840[14]), .I2(n767), .I3(n18391), 
            .O(Gain1_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_10 (.CI(n18391), .I0(n840[14]), .I1(n767), .CO(n18392));
    SB_LUT4 add_1225_9_lut (.I0(GND_net), .I1(n839[14]), .I2(n763), .I3(n18390), 
            .O(Gain1_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_9 (.CI(n18390), .I0(n839[14]), .I1(n763), .CO(n18391));
    SB_LUT4 add_1225_8_lut (.I0(GND_net), .I1(n838[14]), .I2(n759), .I3(n18389), 
            .O(Gain1_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_8 (.CI(n18389), .I0(n838[14]), .I1(n759), .CO(n18390));
    SB_LUT4 add_1225_7_lut (.I0(GND_net), .I1(n837[14]), .I2(n755), .I3(n18388), 
            .O(Gain1_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_7 (.CI(n18388), .I0(n837[14]), .I1(n755), .CO(n18389));
    SB_LUT4 add_1225_6_lut (.I0(GND_net), .I1(n836[14]), .I2(n751), .I3(n18387), 
            .O(Gain1_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_6 (.CI(n18387), .I0(n836[14]), .I1(n751), .CO(n18388));
    SB_LUT4 add_1225_5_lut (.I0(GND_net), .I1(n835[14]), .I2(n747), .I3(n18386), 
            .O(Gain1_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_5 (.CI(n18386), .I0(n835[14]), .I1(n747), .CO(n18387));
    SB_LUT4 add_1225_4_lut (.I0(GND_net), .I1(n834[14]), .I2(n743), .I3(n18385), 
            .O(Gain1_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_4 (.CI(n18385), .I0(n834[14]), .I1(n743), .CO(n18386));
    SB_LUT4 add_1225_3_lut (.I0(GND_net), .I1(n833[14]), .I2(n739), .I3(n18384), 
            .O(Gain1_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_3 (.CI(n18384), .I0(n833[14]), .I1(n739), .CO(n18385));
    SB_LUT4 add_1225_2_lut (.I0(GND_net), .I1(n832[14]), .I2(\betaVoltage[15] ), 
            .I3(GND_net), .O(Gain1_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1225_2 (.CI(GND_net), .I0(n832[14]), .I1(\betaVoltage[15] ), 
            .CO(n18384));
    SB_LUT4 Alpha_15__I_0_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n15966), .O(Add1_cast_1[26])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_12 (.CI(n15966), .I0(GND_net), .I1(n1[10]), 
            .CO(n15967));
    SB_LUT4 Alpha_15__I_0_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n15965), .O(Add1_cast_1[25])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_11 (.CI(n15965), .I0(GND_net), .I1(n1[9]), 
            .CO(n15966));
    SB_LUT4 Beta_15__I_0_add_570_3_lut (.I0(GND_net), .I1(n842[2]), .I2(\betaVoltage[9] ), 
            .I3(n15511), .O(n841[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_3 (.CI(n15511), .I0(n842[2]), .I1(\betaVoltage[9] ), 
            .CO(n15512));
    SB_LUT4 Beta_15__I_0_add_570_2_lut (.I0(GND_net), .I1(\betaVoltage[11] ), 
            .I2(\betaVoltage[9] ), .I3(GND_net), .O(n841[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5933_15_lut (.I0(GND_net), .I1(GND_net), .I2(\betaVoltage[14] ), 
            .I3(n17709), .O(n7479[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_15 (.CI(n17709), .I0(GND_net), .I1(\betaVoltage[14] ), 
            .CO(n7494));
    SB_LUT4 add_5933_14_lut (.I0(GND_net), .I1(\betaVoltage[15] ), .I2(\betaVoltage[14] ), 
            .I3(n17708), .O(n7479[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_14 (.CI(n17708), .I0(\betaVoltage[15] ), .I1(\betaVoltage[14] ), 
            .CO(n17709));
    SB_LUT4 add_5933_13_lut (.I0(GND_net), .I1(GND_net), .I2(GND_net), 
            .I3(n17707), .O(n7479[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_9 (.CI(n15604), .I0(n840[8]), .I1(\betaVoltage[7] ), 
            .CO(n15605));
    SB_LUT4 Beta_15__I_0_add_568_8_lut (.I0(GND_net), .I1(n840[7]), .I2(\betaVoltage[7] ), 
            .I3(n15603), .O(n839[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_570_2 (.CI(GND_net), .I0(\betaVoltage[11] ), 
            .I1(\betaVoltage[9] ), .CO(n15511));
    SB_LUT4 Alpha_15__I_0_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n15964), .O(Add1_cast_1[24])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_10 (.CI(n15964), .I0(GND_net), .I1(n1[8]), 
            .CO(n15965));
    SB_LUT4 Alpha_15__I_0_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n15963), .O(Add1_cast_1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_9 (.CI(n15963), .I0(GND_net), .I1(n1[7]), 
            .CO(n15964));
    SB_LUT4 Beta_15__I_0_add_571_14_lut (.I0(GND_net), .I1(n843[13]), .I2(GND_net), 
            .I3(n15509), .O(n842[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Alpha_15__I_0_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n15962), .O(Add1_cast_1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_8 (.CI(n15962), .I0(GND_net), .I1(n1[6]), 
            .CO(n15963));
    SB_LUT4 Alpha_15__I_0_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n15961), .O(Add1_cast_1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_565_12_lut (.I0(GND_net), .I1(n837[11]), .I2(\betaVoltage[4] ), 
            .I3(n15827), .O(n836[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_14 (.CI(n15509), .I0(n843[13]), .I1(GND_net), 
            .CO(n779));
    SB_CARRY Alpha_15__I_0_add_3_7 (.CI(n15961), .I0(GND_net), .I1(n1[5]), 
            .CO(n15962));
    SB_LUT4 Alpha_15__I_0_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n15960), .O(Add1_cast_1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_13_lut (.I0(GND_net), .I1(n843[12]), .I2(\betaVoltage[10] ), 
            .I3(n15508), .O(n842[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_13 (.CI(n15508), .I0(n843[12]), .I1(\betaVoltage[10] ), 
            .CO(n15509));
    SB_CARRY Alpha_15__I_0_add_3_6 (.CI(n15960), .I0(GND_net), .I1(n1[4]), 
            .CO(n15961));
    SB_LUT4 Alpha_15__I_0_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n15959), .O(Add1_cast_1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_571_12_lut (.I0(GND_net), .I1(n843[11]), .I2(\betaVoltage[10] ), 
            .I3(n15507), .O(n842[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_12 (.CI(n15507), .I0(n843[11]), .I1(\betaVoltage[10] ), 
            .CO(n15508));
    SB_CARRY Alpha_15__I_0_add_3_5 (.CI(n15959), .I0(GND_net), .I1(n1[3]), 
            .CO(n15960));
    SB_LUT4 Alpha_15__I_0_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1007[18]), 
            .I3(n15958), .O(Add1_cast_1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_4 (.CI(n15958), .I0(GND_net), .I1(n1_adj_1007[18]), 
            .CO(n15959));
    SB_LUT4 Alpha_15__I_0_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1007[17]), 
            .I3(n15957), .O(Add1_cast_1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_3 (.CI(n15957), .I0(GND_net), .I1(n1_adj_1007[17]), 
            .CO(n15958));
    SB_LUT4 Alpha_15__I_0_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(Add1_cast_1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam Alpha_15__I_0_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Alpha_15__I_0_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n15957));
    SB_LUT4 Beta_15__I_0_add_571_11_lut (.I0(GND_net), .I1(n843[10]), .I2(GND_net), 
            .I3(n15506), .O(n842[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_12 (.CI(n15827), .I0(n837[11]), .I1(\betaVoltage[4] ), 
            .CO(n15828));
    SB_CARRY Beta_15__I_0_add_571_11 (.CI(n15506), .I0(n843[10]), .I1(GND_net), 
            .CO(n15507));
    SB_LUT4 Beta_15__I_0_add_571_10_lut (.I0(GND_net), .I1(n843[9]), .I2(\betaVoltage[10] ), 
            .I3(n15505), .O(n842[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_10 (.CI(n15505), .I0(n843[9]), .I1(\betaVoltage[10] ), 
            .CO(n15506));
    SB_LUT4 Beta_15__I_0_add_571_9_lut (.I0(GND_net), .I1(n843[8]), .I2(\betaVoltage[10] ), 
            .I3(n15504), .O(n842[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_9 (.CI(n15504), .I0(n843[8]), .I1(\betaVoltage[10] ), 
            .CO(n15505));
    SB_LUT4 Beta_15__I_0_add_571_8_lut (.I0(GND_net), .I1(n843[7]), .I2(\betaVoltage[10] ), 
            .I3(n15503), .O(n842[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_8 (.CI(n15503), .I0(n843[7]), .I1(\betaVoltage[10] ), 
            .CO(n15504));
    SB_LUT4 Beta_15__I_0_add_571_7_lut (.I0(GND_net), .I1(n843[6]), .I2(GND_net), 
            .I3(n15502), .O(n842[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_7 (.CI(n15502), .I0(n843[6]), .I1(GND_net), 
            .CO(n15503));
    SB_LUT4 Beta_15__I_0_add_571_6_lut (.I0(GND_net), .I1(n843[5]), .I2(\betaVoltage[10] ), 
            .I3(n15501), .O(n842[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_6 (.CI(n15501), .I0(n843[5]), .I1(\betaVoltage[10] ), 
            .CO(n15502));
    SB_LUT4 Beta_15__I_0_add_571_5_lut (.I0(GND_net), .I1(n843[4]), .I2(\betaVoltage[10] ), 
            .I3(n15500), .O(n842[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_5 (.CI(n15500), .I0(n843[4]), .I1(\betaVoltage[10] ), 
            .CO(n15501));
    SB_LUT4 Beta_15__I_0_add_571_4_lut (.I0(GND_net), .I1(n843[3]), .I2(GND_net), 
            .I3(n15499), .O(n842[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_4 (.CI(n15499), .I0(n843[3]), .I1(GND_net), 
            .CO(n15500));
    SB_LUT4 Beta_15__I_0_add_571_3_lut (.I0(GND_net), .I1(n843[2]), .I2(\betaVoltage[10] ), 
            .I3(n15498), .O(n842[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_3 (.CI(n15498), .I0(n843[2]), .I1(\betaVoltage[10] ), 
            .CO(n15499));
    SB_LUT4 Beta_15__I_0_add_571_2_lut (.I0(GND_net), .I1(\betaVoltage[12] ), 
            .I2(\betaVoltage[10] ), .I3(GND_net), .O(n842[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_571_2 (.CI(GND_net), .I0(\betaVoltage[12] ), 
            .I1(\betaVoltage[10] ), .CO(n15498));
    SB_LUT4 Beta_15__I_0_add_572_14_lut (.I0(GND_net), .I1(n844[13]), .I2(GND_net), 
            .I3(n15496), .O(n843[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_14 (.CI(n15496), .I0(n844[13]), .I1(GND_net), 
            .CO(n783));
    SB_LUT4 Beta_15__I_0_add_572_13_lut (.I0(GND_net), .I1(n844[12]), .I2(\betaVoltage[11] ), 
            .I3(n15495), .O(n843[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_13 (.CI(n15495), .I0(n844[12]), .I1(\betaVoltage[11] ), 
            .CO(n15496));
    SB_LUT4 Beta_15__I_0_add_572_12_lut (.I0(GND_net), .I1(n844[11]), .I2(\betaVoltage[11] ), 
            .I3(n15494), .O(n843[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_12 (.CI(n15494), .I0(n844[11]), .I1(\betaVoltage[11] ), 
            .CO(n15495));
    SB_LUT4 Beta_15__I_0_add_572_11_lut (.I0(GND_net), .I1(n844[10]), .I2(GND_net), 
            .I3(n15493), .O(n843[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_11 (.CI(n15493), .I0(n844[10]), .I1(GND_net), 
            .CO(n15494));
    SB_LUT4 Beta_15__I_0_add_572_10_lut (.I0(GND_net), .I1(n844[9]), .I2(\betaVoltage[11] ), 
            .I3(n15492), .O(n843[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_10 (.CI(n15492), .I0(n844[9]), .I1(\betaVoltage[11] ), 
            .CO(n15493));
    SB_LUT4 Beta_15__I_0_add_572_9_lut (.I0(GND_net), .I1(n844[8]), .I2(\betaVoltage[11] ), 
            .I3(n15491), .O(n843[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_9 (.CI(n15491), .I0(n844[8]), .I1(\betaVoltage[11] ), 
            .CO(n15492));
    SB_LUT4 Beta_15__I_0_add_572_8_lut (.I0(GND_net), .I1(n844[7]), .I2(\betaVoltage[11] ), 
            .I3(n15490), .O(n843[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_8 (.CI(n15490), .I0(n844[7]), .I1(\betaVoltage[11] ), 
            .CO(n15491));
    SB_LUT4 Beta_15__I_0_add_572_7_lut (.I0(GND_net), .I1(n844[6]), .I2(GND_net), 
            .I3(n15489), .O(n843[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_7 (.CI(n15489), .I0(n844[6]), .I1(GND_net), 
            .CO(n15490));
    SB_LUT4 Beta_15__I_0_add_572_6_lut (.I0(GND_net), .I1(n844[5]), .I2(\betaVoltage[11] ), 
            .I3(n15488), .O(n843[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_565_11_lut (.I0(GND_net), .I1(n837[10]), .I2(GND_net), 
            .I3(n15826), .O(n836[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_6 (.CI(n15488), .I0(n844[5]), .I1(\betaVoltage[11] ), 
            .CO(n15489));
    SB_LUT4 Beta_15__I_0_add_572_5_lut (.I0(GND_net), .I1(n844[4]), .I2(\betaVoltage[11] ), 
            .I3(n15487), .O(n843[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_5 (.CI(n15487), .I0(n844[4]), .I1(\betaVoltage[11] ), 
            .CO(n15488));
    SB_LUT4 Beta_15__I_0_add_572_4_lut (.I0(GND_net), .I1(n844[3]), .I2(GND_net), 
            .I3(n15486), .O(n843[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_4 (.CI(n15486), .I0(n844[3]), .I1(GND_net), 
            .CO(n15487));
    SB_LUT4 Beta_15__I_0_add_572_3_lut (.I0(GND_net), .I1(n844[2]), .I2(\betaVoltage[11] ), 
            .I3(n15485), .O(n843[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_3 (.CI(n15485), .I0(n844[2]), .I1(\betaVoltage[11] ), 
            .CO(n15486));
    SB_LUT4 Beta_15__I_0_add_572_2_lut (.I0(GND_net), .I1(\betaVoltage[13] ), 
            .I2(\betaVoltage[11] ), .I3(GND_net), .O(n843[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_572_2 (.CI(GND_net), .I0(\betaVoltage[13] ), 
            .I1(\betaVoltage[11] ), .CO(n15485));
    SB_LUT4 Beta_15__I_0_add_573_14_lut (.I0(GND_net), .I1(n845[13]), .I2(GND_net), 
            .I3(n15483), .O(n844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_14 (.CI(n15483), .I0(n845[13]), .I1(GND_net), 
            .CO(n787));
    SB_LUT4 Beta_15__I_0_add_573_13_lut (.I0(GND_net), .I1(n845[12]), .I2(\betaVoltage[12] ), 
            .I3(n15482), .O(n844[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_573_13 (.CI(n15482), .I0(n845[12]), .I1(\betaVoltage[12] ), 
            .CO(n15483));
    SB_LUT4 Beta_15__I_0_add_561_14_lut (.I0(GND_net), .I1(n833[13]), .I2(GND_net), 
            .I3(n15881), .O(n832[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_14 (.CI(n15881), .I0(n833[13]), .I1(GND_net), 
            .CO(n739));
    SB_LUT4 Beta_15__I_0_add_561_13_lut (.I0(GND_net), .I1(n833[12]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15880), .O(Gain1_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_13 (.CI(n15880), .I0(n833[12]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15881));
    SB_LUT4 Beta_15__I_0_add_561_12_lut (.I0(GND_net), .I1(n833[11]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15879), .O(\Gain1_mul_temp[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_12 (.CI(n15879), .I0(n833[11]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15880));
    SB_LUT4 Beta_15__I_0_add_561_11_lut (.I0(GND_net), .I1(n833[10]), .I2(GND_net), 
            .I3(n15878), .O(\Gain1_mul_temp[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_11 (.CI(n15878), .I0(n833[10]), .I1(GND_net), 
            .CO(n15879));
    SB_LUT4 Beta_15__I_0_add_561_10_lut (.I0(GND_net), .I1(n833[9]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15877), .O(\Gain1_mul_temp[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_10 (.CI(n15877), .I0(n833[9]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15878));
    SB_LUT4 Beta_15__I_0_add_561_9_lut (.I0(GND_net), .I1(n833[8]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15876), .O(\Gain1_mul_temp[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_9 (.CI(n15876), .I0(n833[8]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15877));
    SB_LUT4 Beta_15__I_0_add_561_8_lut (.I0(GND_net), .I1(n833[7]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15875), .O(\Gain1_mul_temp[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_8 (.CI(n15875), .I0(n833[7]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15876));
    SB_LUT4 Beta_15__I_0_add_561_7_lut (.I0(GND_net), .I1(n833[6]), .I2(GND_net), 
            .I3(n15874), .O(\Gain1_mul_temp[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_7 (.CI(n15874), .I0(n833[6]), .I1(GND_net), 
            .CO(n15875));
    SB_LUT4 Beta_15__I_0_add_561_6_lut (.I0(GND_net), .I1(n833[5]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15873), .O(\Gain1_mul_temp[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_6 (.CI(n15873), .I0(n833[5]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15874));
    SB_LUT4 Beta_15__I_0_add_561_5_lut (.I0(GND_net), .I1(n833[4]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15872), .O(\Gain1_mul_temp[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_5 (.CI(n15872), .I0(n833[4]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15873));
    SB_LUT4 Beta_15__I_0_add_561_4_lut (.I0(GND_net), .I1(n833[3]), .I2(GND_net), 
            .I3(n15871), .O(\Gain1_mul_temp[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_4 (.CI(n15871), .I0(n833[3]), .I1(GND_net), 
            .CO(n15872));
    SB_LUT4 Beta_15__I_0_add_561_3_lut (.I0(GND_net), .I1(n833[2]), .I2(\Gain1_mul_temp[1] ), 
            .I3(n15870), .O(\Gain1_mul_temp[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_3 (.CI(n15870), .I0(n833[2]), .I1(\Gain1_mul_temp[1] ), 
            .CO(n15871));
    SB_LUT4 Beta_15__I_0_add_561_2_lut (.I0(GND_net), .I1(\betaVoltage[2] ), 
            .I2(\Gain1_mul_temp[1] ), .I3(GND_net), .O(\Gain1_mul_temp[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_561_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_561_2 (.CI(GND_net), .I0(\betaVoltage[2] ), 
            .I1(\Gain1_mul_temp[1] ), .CO(n15870));
    SB_LUT4 Beta_15__I_0_add_562_14_lut (.I0(GND_net), .I1(n834[13]), .I2(GND_net), 
            .I3(n15868), .O(n833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_14 (.CI(n15868), .I0(n834[13]), .I1(GND_net), 
            .CO(n743));
    SB_LUT4 Beta_15__I_0_add_562_13_lut (.I0(GND_net), .I1(n834[12]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15867), .O(n833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_13 (.CI(n15867), .I0(n834[12]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15868));
    SB_LUT4 Beta_15__I_0_add_562_12_lut (.I0(GND_net), .I1(n834[11]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15866), .O(n833[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_12 (.CI(n15866), .I0(n834[11]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15867));
    SB_LUT4 Beta_15__I_0_add_562_11_lut (.I0(GND_net), .I1(n834[10]), .I2(GND_net), 
            .I3(n15865), .O(n833[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_11 (.CI(n15865), .I0(n834[10]), .I1(GND_net), 
            .CO(n15866));
    SB_LUT4 Beta_15__I_0_add_562_10_lut (.I0(GND_net), .I1(n834[9]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15864), .O(n833[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_10 (.CI(n15864), .I0(n834[9]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15865));
    SB_LUT4 Beta_15__I_0_add_562_9_lut (.I0(GND_net), .I1(n834[8]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15863), .O(n833[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_9 (.CI(n15863), .I0(n834[8]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15864));
    SB_LUT4 Beta_15__I_0_add_562_8_lut (.I0(GND_net), .I1(n834[7]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15862), .O(n833[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_8 (.CI(n15862), .I0(n834[7]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15863));
    SB_LUT4 Beta_15__I_0_add_562_7_lut (.I0(GND_net), .I1(n834[6]), .I2(GND_net), 
            .I3(n15861), .O(n833[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_7 (.CI(n15861), .I0(n834[6]), .I1(GND_net), 
            .CO(n15862));
    SB_LUT4 Beta_15__I_0_add_562_6_lut (.I0(GND_net), .I1(n834[5]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15860), .O(n833[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_6 (.CI(n15860), .I0(n834[5]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15861));
    SB_LUT4 Beta_15__I_0_add_562_5_lut (.I0(GND_net), .I1(n834[4]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15859), .O(n833[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_5 (.CI(n15859), .I0(n834[4]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15860));
    SB_LUT4 Beta_15__I_0_add_562_4_lut (.I0(GND_net), .I1(n834[3]), .I2(GND_net), 
            .I3(n15858), .O(n833[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_4 (.CI(n15858), .I0(n834[3]), .I1(GND_net), 
            .CO(n15859));
    SB_LUT4 Beta_15__I_0_add_562_3_lut (.I0(GND_net), .I1(n834[2]), .I2(\Gain1_mul_temp[2] ), 
            .I3(n15857), .O(n833[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_3 (.CI(n15857), .I0(n834[2]), .I1(\Gain1_mul_temp[2] ), 
            .CO(n15858));
    SB_LUT4 Beta_15__I_0_add_562_2_lut (.I0(GND_net), .I1(\betaVoltage[3] ), 
            .I2(\Gain1_mul_temp[2] ), .I3(GND_net), .O(n833[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_562_2 (.CI(GND_net), .I0(\betaVoltage[3] ), 
            .I1(\Gain1_mul_temp[2] ), .CO(n15857));
    SB_LUT4 Beta_15__I_0_add_563_14_lut (.I0(GND_net), .I1(n835[13]), .I2(GND_net), 
            .I3(n15855), .O(n834[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_14 (.CI(n15855), .I0(n835[13]), .I1(GND_net), 
            .CO(n747));
    SB_LUT4 Beta_15__I_0_add_563_13_lut (.I0(GND_net), .I1(n835[12]), .I2(\betaVoltage[2] ), 
            .I3(n15854), .O(n834[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_13 (.CI(n15854), .I0(n835[12]), .I1(\betaVoltage[2] ), 
            .CO(n15855));
    SB_LUT4 Beta_15__I_0_add_563_12_lut (.I0(GND_net), .I1(n835[11]), .I2(\betaVoltage[2] ), 
            .I3(n15853), .O(n834[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_12 (.CI(n15853), .I0(n835[11]), .I1(\betaVoltage[2] ), 
            .CO(n15854));
    SB_LUT4 Beta_15__I_0_add_563_11_lut (.I0(GND_net), .I1(n835[10]), .I2(GND_net), 
            .I3(n15852), .O(n834[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_11 (.CI(n15852), .I0(n835[10]), .I1(GND_net), 
            .CO(n15853));
    SB_LUT4 Beta_15__I_0_add_563_10_lut (.I0(GND_net), .I1(n835[9]), .I2(\betaVoltage[2] ), 
            .I3(n15851), .O(n834[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_10 (.CI(n15851), .I0(n835[9]), .I1(\betaVoltage[2] ), 
            .CO(n15852));
    SB_LUT4 Beta_15__I_0_add_563_9_lut (.I0(GND_net), .I1(n835[8]), .I2(\betaVoltage[2] ), 
            .I3(n15850), .O(n834[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_9 (.CI(n15850), .I0(n835[8]), .I1(\betaVoltage[2] ), 
            .CO(n15851));
    SB_LUT4 Beta_15__I_0_add_563_8_lut (.I0(GND_net), .I1(n835[7]), .I2(\betaVoltage[2] ), 
            .I3(n15849), .O(n834[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_8 (.CI(n15849), .I0(n835[7]), .I1(\betaVoltage[2] ), 
            .CO(n15850));
    SB_LUT4 Beta_15__I_0_add_563_7_lut (.I0(GND_net), .I1(n835[6]), .I2(GND_net), 
            .I3(n15848), .O(n834[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_7 (.CI(n15848), .I0(n835[6]), .I1(GND_net), 
            .CO(n15849));
    SB_LUT4 Beta_15__I_0_add_563_6_lut (.I0(GND_net), .I1(n835[5]), .I2(\betaVoltage[2] ), 
            .I3(n15847), .O(n834[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_6 (.CI(n15847), .I0(n835[5]), .I1(\betaVoltage[2] ), 
            .CO(n15848));
    SB_LUT4 Beta_15__I_0_add_563_5_lut (.I0(GND_net), .I1(n835[4]), .I2(\betaVoltage[2] ), 
            .I3(n15846), .O(n834[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_5 (.CI(n15846), .I0(n835[4]), .I1(\betaVoltage[2] ), 
            .CO(n15847));
    SB_LUT4 Beta_15__I_0_add_563_4_lut (.I0(GND_net), .I1(n835[3]), .I2(GND_net), 
            .I3(n15845), .O(n834[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_4 (.CI(n15845), .I0(n835[3]), .I1(GND_net), 
            .CO(n15846));
    SB_LUT4 Beta_15__I_0_add_563_3_lut (.I0(GND_net), .I1(n835[2]), .I2(\betaVoltage[2] ), 
            .I3(n15844), .O(n834[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_3 (.CI(n15844), .I0(n835[2]), .I1(\betaVoltage[2] ), 
            .CO(n15845));
    SB_LUT4 Beta_15__I_0_add_563_2_lut (.I0(GND_net), .I1(\betaVoltage[4] ), 
            .I2(\betaVoltage[2] ), .I3(GND_net), .O(n834[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_563_2 (.CI(GND_net), .I0(\betaVoltage[4] ), 
            .I1(\betaVoltage[2] ), .CO(n15844));
    SB_LUT4 Beta_15__I_0_add_564_14_lut (.I0(GND_net), .I1(n836[13]), .I2(GND_net), 
            .I3(n15842), .O(n835[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_14 (.CI(n15842), .I0(n836[13]), .I1(GND_net), 
            .CO(n751));
    SB_LUT4 Beta_15__I_0_add_564_13_lut (.I0(GND_net), .I1(n836[12]), .I2(\betaVoltage[3] ), 
            .I3(n15841), .O(n835[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_13 (.CI(n15841), .I0(n836[12]), .I1(\betaVoltage[3] ), 
            .CO(n15842));
    SB_LUT4 Beta_15__I_0_add_564_12_lut (.I0(GND_net), .I1(n836[11]), .I2(\betaVoltage[3] ), 
            .I3(n15840), .O(n835[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_12 (.CI(n15840), .I0(n836[11]), .I1(\betaVoltage[3] ), 
            .CO(n15841));
    SB_LUT4 Beta_15__I_0_add_564_11_lut (.I0(GND_net), .I1(n836[10]), .I2(GND_net), 
            .I3(n15839), .O(n835[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_11 (.CI(n15839), .I0(n836[10]), .I1(GND_net), 
            .CO(n15840));
    SB_LUT4 Beta_15__I_0_add_564_10_lut (.I0(GND_net), .I1(n836[9]), .I2(\betaVoltage[3] ), 
            .I3(n15838), .O(n835[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_10 (.CI(n15838), .I0(n836[9]), .I1(\betaVoltage[3] ), 
            .CO(n15839));
    SB_CARRY Beta_15__I_0_add_565_11 (.CI(n15826), .I0(n837[10]), .I1(GND_net), 
            .CO(n15827));
    SB_LUT4 Beta_15__I_0_add_565_10_lut (.I0(GND_net), .I1(n837[9]), .I2(\betaVoltage[4] ), 
            .I3(n15825), .O(n836[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_10 (.CI(n15825), .I0(n837[9]), .I1(\betaVoltage[4] ), 
            .CO(n15826));
    SB_LUT4 Beta_15__I_0_add_565_9_lut (.I0(GND_net), .I1(n837[8]), .I2(\betaVoltage[4] ), 
            .I3(n15824), .O(n836[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_9 (.CI(n15824), .I0(n837[8]), .I1(\betaVoltage[4] ), 
            .CO(n15825));
    SB_LUT4 Beta_15__I_0_add_565_8_lut (.I0(GND_net), .I1(n837[7]), .I2(\betaVoltage[4] ), 
            .I3(n15823), .O(n836[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_8 (.CI(n15823), .I0(n837[7]), .I1(\betaVoltage[4] ), 
            .CO(n15824));
    SB_LUT4 Beta_15__I_0_add_565_7_lut (.I0(GND_net), .I1(n837[6]), .I2(GND_net), 
            .I3(n15822), .O(n836[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_7 (.CI(n15822), .I0(n837[6]), .I1(GND_net), 
            .CO(n15823));
    SB_LUT4 Beta_15__I_0_add_565_6_lut (.I0(GND_net), .I1(n837[5]), .I2(\betaVoltage[4] ), 
            .I3(n15821), .O(n836[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_6 (.CI(n15821), .I0(n837[5]), .I1(\betaVoltage[4] ), 
            .CO(n15822));
    SB_LUT4 Beta_15__I_0_add_565_5_lut (.I0(GND_net), .I1(n837[4]), .I2(\betaVoltage[4] ), 
            .I3(n15820), .O(n836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_5 (.CI(n15820), .I0(n837[4]), .I1(\betaVoltage[4] ), 
            .CO(n15821));
    SB_LUT4 Beta_15__I_0_add_564_6_lut (.I0(GND_net), .I1(n836[5]), .I2(\betaVoltage[3] ), 
            .I3(n15834), .O(n835[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_13 (.CI(n17707), .I0(GND_net), .I1(GND_net), .CO(n17708));
    SB_LUT4 add_5933_12_lut (.I0(GND_net), .I1(GND_net), .I2(\betaVoltage[14] ), 
            .I3(n17706), .O(n7479[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_12 (.CI(n17706), .I0(GND_net), .I1(\betaVoltage[14] ), 
            .CO(n17707));
    SB_LUT4 add_5933_11_lut (.I0(GND_net), .I1(GND_net), .I2(\betaVoltage[14] ), 
            .I3(n17705), .O(n7479[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_11 (.CI(n17705), .I0(GND_net), .I1(\betaVoltage[14] ), 
            .CO(n17706));
    SB_LUT4 add_5933_10_lut (.I0(GND_net), .I1(\betaVoltage[15] ), .I2(\betaVoltage[14] ), 
            .I3(n17704), .O(n7479[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5933_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5933_10 (.CI(n17704), .I0(\betaVoltage[15] ), .I1(\betaVoltage[14] ), 
            .CO(n17705));
    SB_LUT4 Beta_15__I_0_add_565_4_lut (.I0(GND_net), .I1(n837[3]), .I2(GND_net), 
            .I3(n15819), .O(n836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_4 (.CI(n15819), .I0(n837[3]), .I1(GND_net), 
            .CO(n15820));
    SB_LUT4 Beta_15__I_0_add_565_3_lut (.I0(GND_net), .I1(n837[2]), .I2(\betaVoltage[4] ), 
            .I3(n15818), .O(n836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_3 (.CI(n15818), .I0(n837[2]), .I1(\betaVoltage[4] ), 
            .CO(n15819));
    SB_LUT4 Beta_15__I_0_add_565_2_lut (.I0(GND_net), .I1(\betaVoltage[6] ), 
            .I2(\betaVoltage[4] ), .I3(GND_net), .O(n836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_565_2 (.CI(GND_net), .I0(\betaVoltage[6] ), 
            .I1(\betaVoltage[4] ), .CO(n15818));
    SB_LUT4 Beta_15__I_0_add_566_14_lut (.I0(GND_net), .I1(n838[13]), .I2(GND_net), 
            .I3(n15816), .O(n837[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_14 (.CI(n15816), .I0(n838[13]), .I1(GND_net), 
            .CO(n759));
    SB_LUT4 Beta_15__I_0_add_566_13_lut (.I0(GND_net), .I1(n838[12]), .I2(\betaVoltage[5] ), 
            .I3(n15815), .O(n837[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_13 (.CI(n15815), .I0(n838[12]), .I1(\betaVoltage[5] ), 
            .CO(n15816));
    SB_LUT4 Beta_15__I_0_add_566_12_lut (.I0(GND_net), .I1(n838[11]), .I2(\betaVoltage[5] ), 
            .I3(n15814), .O(n837[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_12 (.CI(n15814), .I0(n838[11]), .I1(\betaVoltage[5] ), 
            .CO(n15815));
    SB_LUT4 Beta_15__I_0_add_566_11_lut (.I0(GND_net), .I1(n838[10]), .I2(GND_net), 
            .I3(n15813), .O(n837[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_11 (.CI(n15813), .I0(n838[10]), .I1(GND_net), 
            .CO(n15814));
    SB_LUT4 Beta_15__I_0_add_566_10_lut (.I0(GND_net), .I1(n838[9]), .I2(\betaVoltage[5] ), 
            .I3(n15812), .O(n837[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_10 (.CI(n15812), .I0(n838[9]), .I1(\betaVoltage[5] ), 
            .CO(n15813));
    SB_LUT4 Beta_15__I_0_add_566_9_lut (.I0(GND_net), .I1(n838[8]), .I2(\betaVoltage[5] ), 
            .I3(n15811), .O(n837[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_9 (.CI(n15811), .I0(n838[8]), .I1(\betaVoltage[5] ), 
            .CO(n15812));
    SB_LUT4 Beta_15__I_0_add_566_8_lut (.I0(GND_net), .I1(n838[7]), .I2(\betaVoltage[5] ), 
            .I3(n15810), .O(n837[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_8 (.CI(n15810), .I0(n838[7]), .I1(\betaVoltage[5] ), 
            .CO(n15811));
    SB_LUT4 Beta_15__I_0_add_566_7_lut (.I0(GND_net), .I1(n838[6]), .I2(GND_net), 
            .I3(n15809), .O(n837[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_7 (.CI(n15809), .I0(n838[6]), .I1(GND_net), 
            .CO(n15810));
    SB_LUT4 Beta_15__I_0_add_566_6_lut (.I0(GND_net), .I1(n838[5]), .I2(\betaVoltage[5] ), 
            .I3(n15808), .O(n837[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_6 (.CI(n15808), .I0(n838[5]), .I1(\betaVoltage[5] ), 
            .CO(n15809));
    SB_LUT4 Beta_15__I_0_add_566_5_lut (.I0(GND_net), .I1(n838[4]), .I2(\betaVoltage[5] ), 
            .I3(n15807), .O(n837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_9_lut (.I0(GND_net), .I1(n836[8]), .I2(\betaVoltage[3] ), 
            .I3(n15837), .O(n835[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_5 (.CI(n15807), .I0(n838[4]), .I1(\betaVoltage[5] ), 
            .CO(n15808));
    SB_LUT4 Beta_15__I_0_add_566_4_lut (.I0(GND_net), .I1(n838[3]), .I2(GND_net), 
            .I3(n15806), .O(n837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_4 (.CI(n15806), .I0(n838[3]), .I1(GND_net), 
            .CO(n15807));
    SB_LUT4 Beta_15__I_0_add_566_3_lut (.I0(GND_net), .I1(n838[2]), .I2(\betaVoltage[5] ), 
            .I3(n15805), .O(n837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_3 (.CI(n15805), .I0(n838[2]), .I1(\betaVoltage[5] ), 
            .CO(n15806));
    SB_LUT4 Beta_15__I_0_add_566_2_lut (.I0(GND_net), .I1(\betaVoltage[7] ), 
            .I2(\betaVoltage[5] ), .I3(GND_net), .O(n837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_566_2 (.CI(GND_net), .I0(\betaVoltage[7] ), 
            .I1(\betaVoltage[5] ), .CO(n15805));
    SB_LUT4 Beta_15__I_0_add_564_8_lut (.I0(GND_net), .I1(n836[7]), .I2(\betaVoltage[3] ), 
            .I3(n15836), .O(n835[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_8 (.CI(n15836), .I0(n836[7]), .I1(\betaVoltage[3] ), 
            .CO(n15837));
    SB_LUT4 Beta_15__I_0_add_564_7_lut (.I0(GND_net), .I1(n836[6]), .I2(GND_net), 
            .I3(n15835), .O(n835[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_7 (.CI(n15835), .I0(n836[6]), .I1(GND_net), 
            .CO(n15836));
    SB_LUT4 sub_67_add_2_19_lut (.I0(GND_net), .I1(Gain1_mul_temp[30]), 
            .I2(n1[15]), .I3(n15719), .O(\abcVoltage_1[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_18_lut (.I0(GND_net), .I1(Gain1_mul_temp[30]), 
            .I2(n1[15]), .I3(n15718), .O(\abcVoltage_1[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_18 (.CI(n15718), .I0(Gain1_mul_temp[30]), .I1(n1[15]), 
            .CO(n15719));
    SB_LUT4 sub_67_add_2_17_lut (.I0(GND_net), .I1(Gain1_mul_temp[29]), 
            .I2(n1[15]), .I3(n15717), .O(\abcVoltage_1[29] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_17 (.CI(n15717), .I0(Gain1_mul_temp[29]), .I1(n1[15]), 
            .CO(n15718));
    SB_LUT4 sub_67_add_2_16_lut (.I0(GND_net), .I1(Gain1_mul_temp[28]), 
            .I2(n1[14]), .I3(n15716), .O(\abcVoltage_1[28] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_16 (.CI(n15716), .I0(Gain1_mul_temp[28]), .I1(n1[14]), 
            .CO(n15717));
    SB_CARRY Beta_15__I_0_add_568_12 (.CI(n15607), .I0(n840[11]), .I1(\betaVoltage[7] ), 
            .CO(n15608));
    SB_LUT4 sub_67_add_2_15_lut (.I0(GND_net), .I1(Gain1_mul_temp[27]), 
            .I2(n1[13]), .I3(n15715), .O(\abcVoltage_1[27] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_15 (.CI(n15715), .I0(Gain1_mul_temp[27]), .I1(n1[13]), 
            .CO(n15716));
    SB_LUT4 sub_67_add_2_14_lut (.I0(GND_net), .I1(Gain1_mul_temp[26]), 
            .I2(n1[12]), .I3(n15714), .O(\abcVoltage_1[26] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_14 (.CI(n15714), .I0(Gain1_mul_temp[26]), .I1(n1[12]), 
            .CO(n15715));
    SB_LUT4 sub_67_add_2_13_lut (.I0(GND_net), .I1(Gain1_mul_temp[25]), 
            .I2(n1[11]), .I3(n15713), .O(\abcVoltage_1[25] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_13 (.CI(n15713), .I0(Gain1_mul_temp[25]), .I1(n1[11]), 
            .CO(n15714));
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(Gain1_mul_temp[24]), 
            .I2(n1[10]), .I3(n15712), .O(\abcVoltage_1[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_12 (.CI(n15712), .I0(Gain1_mul_temp[24]), .I1(n1[10]), 
            .CO(n15713));
    SB_LUT4 sub_67_add_2_11_lut (.I0(GND_net), .I1(Gain1_mul_temp[23]), 
            .I2(n1[9]), .I3(n15711), .O(\abcVoltage_1[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_11 (.CI(n15711), .I0(Gain1_mul_temp[23]), .I1(n1[9]), 
            .CO(n15712));
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(Gain1_mul_temp[22]), 
            .I2(n1[8]), .I3(n15710), .O(\abcVoltage_1[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n15710), .I0(Gain1_mul_temp[22]), .I1(n1[8]), 
            .CO(n15711));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(Gain1_mul_temp[21]), .I2(n1[7]), 
            .I3(n15709), .O(\abcVoltage_1[21] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n15709), .I0(Gain1_mul_temp[21]), .I1(n1[7]), 
            .CO(n15710));
    SB_LUT4 sub_67_add_2_8_lut (.I0(GND_net), .I1(Gain1_mul_temp[20]), .I2(n1[6]), 
            .I3(n15708), .O(\abcVoltage_1[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_8 (.CI(n15708), .I0(Gain1_mul_temp[20]), .I1(n1[6]), 
            .CO(n15709));
    SB_LUT4 sub_67_add_2_7_lut (.I0(GND_net), .I1(Gain1_mul_temp[19]), .I2(n1[5]), 
            .I3(n15707), .O(\abcVoltage_1[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_7 (.CI(n15707), .I0(Gain1_mul_temp[19]), .I1(n1[5]), 
            .CO(n15708));
    SB_LUT4 Beta_15__I_0_add_567_14_lut (.I0(GND_net), .I1(n839[13]), .I2(GND_net), 
            .I3(n15622), .O(n838[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_6_lut (.I0(GND_net), .I1(Gain1_mul_temp[18]), .I2(n1[4]), 
            .I3(n15706), .O(\abcVoltage_1[18] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_6 (.CI(n15706), .I0(Gain1_mul_temp[18]), .I1(n1[4]), 
            .CO(n15707));
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(Gain1_mul_temp[17]), .I2(n1[3]), 
            .I3(n15705), .O(\abcVoltage_1[17] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_5 (.CI(n15705), .I0(Gain1_mul_temp[17]), .I1(n1[3]), 
            .CO(n15706));
    SB_CARRY Beta_15__I_0_add_567_14 (.CI(n15622), .I0(n839[13]), .I1(GND_net), 
            .CO(n763));
    SB_LUT4 Beta_15__I_0_add_567_13_lut (.I0(GND_net), .I1(n839[12]), .I2(\betaVoltage[6] ), 
            .I3(n15621), .O(n838[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(Gain1_mul_temp[16]), .I2(n1_adj_1007[18]), 
            .I3(n15704), .O(\abcVoltage_1[16] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_4 (.CI(n15704), .I0(Gain1_mul_temp[16]), .I1(n1_adj_1007[18]), 
            .CO(n15705));
    SB_LUT4 sub_67_add_2_3_lut (.I0(GND_net), .I1(Gain1_mul_temp[15]), .I2(n1_adj_1007[17]), 
            .I3(n15703), .O(\abcVoltage_1[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_3 (.CI(n15703), .I0(Gain1_mul_temp[15]), .I1(n1_adj_1007[17]), 
            .CO(n15704));
    SB_LUT4 sub_67_add_2_2_lut (.I0(GND_net), .I1(Gain1_mul_temp[14]), .I2(n1[0]), 
            .I3(VCC_net), .O(\abcVoltage_1[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(Gain1_mul_temp[14]), .I1(n1[0]), 
            .CO(n15703));
    SB_LUT4 sub_68_add_2_33_lut (.I0(GND_net), .I1(Add1_cast_1[32]), .I2(n1_adj_1008[31]), 
            .I3(n15702), .O(\abcVoltage_2[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_68_add_2_32_lut (.I0(GND_net), .I1(Add1_cast_1[32]), .I2(n1_adj_1008[31]), 
            .I3(n15701), .O(\abcVoltage_2[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_32 (.CI(n15701), .I0(Add1_cast_1[32]), .I1(n1_adj_1008[31]), 
            .CO(n15702));
    SB_LUT4 sub_68_add_2_31_lut (.I0(GND_net), .I1(Add1_cast_1[31]), .I2(n1_adj_1008[29]), 
            .I3(n15700), .O(\abcVoltage_2[29] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_31 (.CI(n15700), .I0(Add1_cast_1[31]), .I1(n1_adj_1008[29]), 
            .CO(n15701));
    SB_LUT4 sub_68_add_2_30_lut (.I0(GND_net), .I1(Add1_cast_1[30]), .I2(n1_adj_1008[28]), 
            .I3(n15699), .O(\abcVoltage_2[28] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_30 (.CI(n15699), .I0(Add1_cast_1[30]), .I1(n1_adj_1008[28]), 
            .CO(n15700));
    SB_LUT4 sub_68_add_2_29_lut (.I0(GND_net), .I1(Add1_cast_1[29]), .I2(n1_adj_1008[27]), 
            .I3(n15698), .O(\abcVoltage_2[27] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_29 (.CI(n15698), .I0(Add1_cast_1[29]), .I1(n1_adj_1008[27]), 
            .CO(n15699));
    SB_LUT4 sub_68_add_2_28_lut (.I0(GND_net), .I1(Add1_cast_1[28]), .I2(n1_adj_1008[26]), 
            .I3(n15697), .O(\abcVoltage_2[26] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_28 (.CI(n15697), .I0(Add1_cast_1[28]), .I1(n1_adj_1008[26]), 
            .CO(n15698));
    SB_LUT4 sub_68_add_2_27_lut (.I0(GND_net), .I1(Add1_cast_1[27]), .I2(n1_adj_1008[25]), 
            .I3(n15696), .O(\abcVoltage_2[25] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_27 (.CI(n15696), .I0(Add1_cast_1[27]), .I1(n1_adj_1008[25]), 
            .CO(n15697));
    SB_LUT4 Beta_15__I_0_add_564_4_lut (.I0(GND_net), .I1(n836[3]), .I2(GND_net), 
            .I3(n15832), .O(n835[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_564_6 (.CI(n15834), .I0(n836[5]), .I1(\betaVoltage[3] ), 
            .CO(n15835));
    SB_LUT4 sub_68_add_2_26_lut (.I0(GND_net), .I1(Add1_cast_1[26]), .I2(n1_adj_1008[24]), 
            .I3(n15695), .O(\abcVoltage_2[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_26 (.CI(n15695), .I0(Add1_cast_1[26]), .I1(n1_adj_1008[24]), 
            .CO(n15696));
    SB_LUT4 sub_68_add_2_25_lut (.I0(GND_net), .I1(Add1_cast_1[25]), .I2(n1_adj_1008[23]), 
            .I3(n15694), .O(\abcVoltage_2[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_25 (.CI(n15694), .I0(Add1_cast_1[25]), .I1(n1_adj_1008[23]), 
            .CO(n15695));
    SB_LUT4 sub_68_add_2_24_lut (.I0(GND_net), .I1(Add1_cast_1[24]), .I2(n1_adj_1008[22]), 
            .I3(n15693), .O(\abcVoltage_2[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_24 (.CI(n15693), .I0(Add1_cast_1[24]), .I1(n1_adj_1008[22]), 
            .CO(n15694));
    SB_LUT4 sub_68_add_2_23_lut (.I0(GND_net), .I1(Add1_cast_1[23]), .I2(n1_adj_1008[21]), 
            .I3(n15692), .O(\abcVoltage_2[21] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_23 (.CI(n15692), .I0(Add1_cast_1[23]), .I1(n1_adj_1008[21]), 
            .CO(n15693));
    SB_LUT4 sub_68_add_2_22_lut (.I0(GND_net), .I1(Add1_cast_1[22]), .I2(n1_adj_1008[20]), 
            .I3(n15691), .O(\abcVoltage_2[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_22 (.CI(n15691), .I0(Add1_cast_1[22]), .I1(n1_adj_1008[20]), 
            .CO(n15692));
    SB_LUT4 sub_68_add_2_21_lut (.I0(GND_net), .I1(Add1_cast_1[21]), .I2(n1_adj_1008[19]), 
            .I3(n15690), .O(\abcVoltage_2[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_21 (.CI(n15690), .I0(Add1_cast_1[21]), .I1(n1_adj_1008[19]), 
            .CO(n15691));
    SB_LUT4 sub_68_add_2_20_lut (.I0(GND_net), .I1(Add1_cast_1[20]), .I2(n1_adj_1008[18]), 
            .I3(n15689), .O(\abcVoltage_2[18] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_20 (.CI(n15689), .I0(Add1_cast_1[20]), .I1(n1_adj_1008[18]), 
            .CO(n15690));
    SB_LUT4 sub_68_add_2_19_lut (.I0(GND_net), .I1(Add1_cast_1[19]), .I2(n1_adj_1008[17]), 
            .I3(n15688), .O(\abcVoltage_2[17] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_19 (.CI(n15688), .I0(Add1_cast_1[19]), .I1(n1_adj_1008[17]), 
            .CO(n15689));
    SB_LUT4 sub_68_add_2_18_lut (.I0(GND_net), .I1(Add1_cast_1[18]), .I2(n1_adj_1008[16]), 
            .I3(n15687), .O(\abcVoltage_2[16] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_18 (.CI(n15687), .I0(Add1_cast_1[18]), .I1(n1_adj_1008[16]), 
            .CO(n15688));
    SB_LUT4 sub_68_add_2_17_lut (.I0(GND_net), .I1(Add1_cast_1[17]), .I2(n1_adj_1008[15]), 
            .I3(n15686), .O(\abcVoltage_2[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_17 (.CI(n15686), .I0(Add1_cast_1[17]), .I1(n1_adj_1008[15]), 
            .CO(n15687));
    SB_LUT4 sub_68_add_2_16_lut (.I0(GND_net), .I1(Add1_cast_1[16]), .I2(n1_adj_1008[14]), 
            .I3(n15685), .O(\abcVoltage_2[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_16 (.CI(n15685), .I0(Add1_cast_1[16]), .I1(n1_adj_1008[14]), 
            .CO(n15686));
    SB_LUT4 sub_68_add_2_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[13]), 
            .I3(n15684), .O(\abcVoltage_2[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_15 (.CI(n15684), .I0(GND_net), .I1(n1_adj_1008[13]), 
            .CO(n15685));
    SB_LUT4 sub_68_add_2_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[12]), 
            .I3(n15683), .O(\abcVoltage_2[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_14 (.CI(n15683), .I0(GND_net), .I1(n1_adj_1008[12]), 
            .CO(n15684));
    SB_LUT4 sub_68_add_2_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[11]), 
            .I3(n15682), .O(\abcVoltage_2[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_13 (.CI(n15682), .I0(GND_net), .I1(n1_adj_1008[11]), 
            .CO(n15683));
    SB_LUT4 sub_68_add_2_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[10]), 
            .I3(n15681), .O(\abcVoltage_2[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_12 (.CI(n15681), .I0(GND_net), .I1(n1_adj_1008[10]), 
            .CO(n15682));
    SB_LUT4 sub_68_add_2_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[9]), 
            .I3(n15680), .O(\abcVoltage_2[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_11 (.CI(n15680), .I0(GND_net), .I1(n1_adj_1008[9]), 
            .CO(n15681));
    SB_LUT4 sub_68_add_2_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[8]), 
            .I3(n15679), .O(\abcVoltage_2[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_10 (.CI(n15679), .I0(GND_net), .I1(n1_adj_1008[8]), 
            .CO(n15680));
    SB_LUT4 sub_68_add_2_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[7]), 
            .I3(n15678), .O(\abcVoltage_2[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_9 (.CI(n15678), .I0(GND_net), .I1(n1_adj_1008[7]), 
            .CO(n15679));
    SB_CARRY Beta_15__I_0_add_564_9 (.CI(n15837), .I0(n836[8]), .I1(\betaVoltage[3] ), 
            .CO(n15838));
    SB_CARRY Beta_15__I_0_add_567_13 (.CI(n15621), .I0(n839[12]), .I1(\betaVoltage[6] ), 
            .CO(n15622));
    SB_LUT4 Beta_15__I_0_add_567_12_lut (.I0(GND_net), .I1(n839[11]), .I2(\betaVoltage[6] ), 
            .I3(n15620), .O(n838[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_12 (.CI(n15620), .I0(n839[11]), .I1(\betaVoltage[6] ), 
            .CO(n15621));
    SB_LUT4 Beta_15__I_0_add_567_11_lut (.I0(GND_net), .I1(n839[10]), .I2(GND_net), 
            .I3(n15619), .O(n838[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_11 (.CI(n15619), .I0(n839[10]), .I1(GND_net), 
            .CO(n15620));
    SB_LUT4 Beta_15__I_0_add_567_10_lut (.I0(GND_net), .I1(n839[9]), .I2(\betaVoltage[6] ), 
            .I3(n15618), .O(n838[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_10 (.CI(n15618), .I0(n839[9]), .I1(\betaVoltage[6] ), 
            .CO(n15619));
    SB_LUT4 Beta_15__I_0_add_567_9_lut (.I0(GND_net), .I1(n839[8]), .I2(\betaVoltage[6] ), 
            .I3(n15617), .O(n838[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_9 (.CI(n15617), .I0(n839[8]), .I1(\betaVoltage[6] ), 
            .CO(n15618));
    SB_LUT4 Beta_15__I_0_add_567_8_lut (.I0(GND_net), .I1(n839[7]), .I2(\betaVoltage[6] ), 
            .I3(n15616), .O(n838[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_68_add_2_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[6]), 
            .I3(n15677), .O(\abcVoltage_2[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_564_5_lut (.I0(GND_net), .I1(n836[4]), .I2(\betaVoltage[3] ), 
            .I3(n15833), .O(n835[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_8 (.CI(n15616), .I0(n839[7]), .I1(\betaVoltage[6] ), 
            .CO(n15617));
    SB_CARRY sub_68_add_2_8 (.CI(n15677), .I0(GND_net), .I1(n1_adj_1008[6]), 
            .CO(n15678));
    SB_LUT4 Beta_15__I_0_add_567_7_lut (.I0(GND_net), .I1(n839[6]), .I2(GND_net), 
            .I3(n15615), .O(n838[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_68_add_2_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[5]), 
            .I3(n15676), .O(\abcVoltage_2[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_568_11_lut (.I0(GND_net), .I1(n840[10]), .I2(GND_net), 
            .I3(n15606), .O(n839[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_7 (.CI(n15615), .I0(n839[6]), .I1(GND_net), 
            .CO(n15616));
    SB_CARRY sub_68_add_2_7 (.CI(n15676), .I0(GND_net), .I1(n1_adj_1008[5]), 
            .CO(n15677));
    SB_LUT4 sub_68_add_2_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[4]), 
            .I3(n15675), .O(\abcVoltage_2[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_6_lut (.I0(GND_net), .I1(n839[5]), .I2(\betaVoltage[6] ), 
            .I3(n15614), .O(n838[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_6 (.CI(n15675), .I0(GND_net), .I1(n1_adj_1008[4]), 
            .CO(n15676));
    SB_LUT4 sub_68_add_2_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[3]), 
            .I3(n15674), .O(\abcVoltage_2[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_6 (.CI(n15614), .I0(n839[5]), .I1(\betaVoltage[6] ), 
            .CO(n15615));
    SB_CARRY sub_68_add_2_5 (.CI(n15674), .I0(GND_net), .I1(n1_adj_1008[3]), 
            .CO(n15675));
    SB_LUT4 sub_68_add_2_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[2]), 
            .I3(n15673), .O(\abcVoltage_2[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Beta_15__I_0_add_567_5_lut (.I0(GND_net), .I1(n839[4]), .I2(\betaVoltage[6] ), 
            .I3(n15613), .O(n838[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_68_add_2_4 (.CI(n15673), .I0(GND_net), .I1(n1_adj_1008[2]), 
            .CO(n15674));
    SB_LUT4 sub_68_add_2_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_1008[1]), 
            .I3(n15672), .O(\abcVoltage_2[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_68_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_5 (.CI(n15613), .I0(n839[4]), .I1(\betaVoltage[6] ), 
            .CO(n15614));
    SB_CARRY sub_68_add_2_3 (.CI(n15672), .I0(GND_net), .I1(n1_adj_1008[1]), 
            .CO(n15673));
    SB_CARRY sub_68_add_2_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), 
            .CO(n15672));
    SB_LUT4 Beta_15__I_0_add_567_4_lut (.I0(GND_net), .I1(n839[3]), .I2(GND_net), 
            .I3(n15612), .O(n838[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_4 (.CI(n15612), .I0(n839[3]), .I1(GND_net), 
            .CO(n15613));
    SB_LUT4 Beta_15__I_0_add_567_3_lut (.I0(GND_net), .I1(n839[2]), .I2(\betaVoltage[6] ), 
            .I3(n15611), .O(n838[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_3 (.CI(n15611), .I0(n839[2]), .I1(\betaVoltage[6] ), 
            .CO(n15612));
    SB_LUT4 Beta_15__I_0_add_567_2_lut (.I0(GND_net), .I1(\betaVoltage[8] ), 
            .I2(\betaVoltage[6] ), .I3(GND_net), .O(n838[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_567_2 (.CI(GND_net), .I0(\betaVoltage[8] ), 
            .I1(\betaVoltage[6] ), .CO(n15611));
    SB_LUT4 Beta_15__I_0_add_568_14_lut (.I0(GND_net), .I1(n840[13]), .I2(GND_net), 
            .I3(n15609), .O(n839[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_14 (.CI(n15609), .I0(n840[13]), .I1(GND_net), 
            .CO(n767));
    SB_CARRY Beta_15__I_0_add_573_2 (.CI(GND_net), .I0(n7479[0]), .I1(\betaVoltage[12] ), 
            .CO(n15472));
    SB_LUT4 Beta_15__I_0_add_568_13_lut (.I0(GND_net), .I1(n840[12]), .I2(\betaVoltage[7] ), 
            .I3(n15608), .O(n839[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_13 (.CI(n15608), .I0(n840[12]), .I1(\betaVoltage[7] ), 
            .CO(n15609));
    SB_LUT4 Beta_15__I_0_add_568_12_lut (.I0(GND_net), .I1(n840[11]), .I2(\betaVoltage[7] ), 
            .I3(n15607), .O(n839[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Beta_15__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Beta_15__I_0_add_568_8 (.CI(n15603), .I0(n840[7]), .I1(\betaVoltage[7] ), 
            .CO(n15604));
    SB_LUT4 sub_68_inv_0_i2_1_lut (.I0(\Gain1_mul_temp[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[1]));
    defparam sub_68_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i3_1_lut (.I0(\Gain1_mul_temp[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[2]));
    defparam sub_68_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i4_1_lut (.I0(\Gain1_mul_temp[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[3]));
    defparam sub_68_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i5_1_lut (.I0(\Gain1_mul_temp[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[4]));
    defparam sub_68_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i6_1_lut (.I0(\Gain1_mul_temp[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[5]));
    defparam sub_68_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i7_1_lut (.I0(\Gain1_mul_temp[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[6]));
    defparam sub_68_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i8_1_lut (.I0(\Gain1_mul_temp[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[7]));
    defparam sub_68_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i9_1_lut (.I0(\Gain1_mul_temp[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[8]));
    defparam sub_68_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i10_1_lut (.I0(\Gain1_mul_temp[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[9]));
    defparam sub_68_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i11_1_lut (.I0(\Gain1_mul_temp[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[10]));
    defparam sub_68_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i12_1_lut (.I0(\Gain1_mul_temp[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[11]));
    defparam sub_68_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i13_1_lut (.I0(\Gain1_mul_temp[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[12]));
    defparam sub_68_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i14_1_lut (.I0(\Gain1_mul_temp[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[13]));
    defparam sub_68_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i15_1_lut (.I0(Gain1_mul_temp[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[14]));
    defparam sub_68_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i16_1_lut (.I0(Gain1_mul_temp[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[15]));
    defparam sub_68_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i17_1_lut (.I0(Gain1_mul_temp[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[16]));
    defparam sub_68_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i18_1_lut (.I0(Gain1_mul_temp[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[17]));
    defparam sub_68_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i19_1_lut (.I0(Gain1_mul_temp[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[18]));
    defparam sub_68_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i20_1_lut (.I0(Gain1_mul_temp[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[19]));
    defparam sub_68_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i21_1_lut (.I0(Gain1_mul_temp[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[20]));
    defparam sub_68_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i22_1_lut (.I0(Gain1_mul_temp[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[21]));
    defparam sub_68_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i23_1_lut (.I0(Gain1_mul_temp[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[22]));
    defparam sub_68_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i24_1_lut (.I0(Gain1_mul_temp[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[23]));
    defparam sub_68_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i25_1_lut (.I0(Gain1_mul_temp[24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[24]));
    defparam sub_68_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i26_1_lut (.I0(Gain1_mul_temp[25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[25]));
    defparam sub_68_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i27_1_lut (.I0(Gain1_mul_temp[26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[26]));
    defparam sub_68_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i28_1_lut (.I0(Gain1_mul_temp[27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[27]));
    defparam sub_68_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i29_1_lut (.I0(Gain1_mul_temp[28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[28]));
    defparam sub_68_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i30_1_lut (.I0(Gain1_mul_temp[29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[29]));
    defparam sub_68_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_68_inv_0_i32_1_lut (.I0(Gain1_mul_temp[30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1008[31]));
    defparam sub_68_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(alphaVoltage[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[0]));
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 Alpha_15__I_0_inv_0_i18_1_lut (.I0(alphaVoltage[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1007[17]));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Clarke_Transform.v(78[25:38])
    defparam Alpha_15__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 Alpha_15__I_0_inv_0_i19_1_lut (.I0(alphaVoltage[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1007[18]));   // ../../hdlcoderFocCurrentFixptHdl/Inverse_Clarke_Transform.v(78[25:38])
    defparam Alpha_15__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(alphaVoltage[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(alphaVoltage[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(alphaVoltage[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(alphaVoltage[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(alphaVoltage[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(alphaVoltage[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(alphaVoltage[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    VCC i1 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module DQ_Current_Control
//

module DQ_Current_Control (GND_net, n14381, pin3_clk_16mhz_N_keep, \Product_mul_temp[26] , 
            \Error_sub_temp[31] , \preSatVoltage[10] , Out_31__N_333, 
            Out_31__N_332, \qVoltage[8] , \qVoltage[5] , \qVoltage[2] , 
            \qVoltage[12] , n14380, \preSatVoltage[23] , \qVoltage[14] , 
            \qVoltage[9] , n14379, \preSatVoltage[13] , \preSatVoltage[12] , 
            \qVoltage[4] , \qVoltage[3] , \qVoltage[15] , n14378, n14377, 
            n14376, n14375, n14374, \qVoltage[6] , n14373, \preSatVoltage[22] , 
            \preSatVoltage[19] , \qVoltage[13] , \qVoltage[10] , \qVoltage[7] , 
            n14354, n14372, n14371, n14370, n14369, n14353, n14368, 
            n14367, n14366, n14365, n14364, n14363, n14362, n14361, 
            n14360, n14359, n14352, n14358, \Amp25_out1[14] , n146, 
            n14357, n14356, n793, n141, n794, \Add_add_temp[34] , 
            \Add_add_temp[33] , \Add_add_temp[32] , \Add_add_temp[31] , 
            \Add_add_temp[30] , \Add_add_temp[29] , \Add_add_temp[28] , 
            \Add_add_temp[27] , \Add_add_temp[26] , \Add_add_temp[25] , 
            \Add_add_temp[24] , \Add_add_temp[23] , \Add_add_temp[22] , 
            \Add_add_temp[21] , \Add_add_temp[20] , \Add_add_temp[19] , 
            \Add_add_temp[18] , \Add_add_temp[17] , \Add_add_temp[16] , 
            \Add_add_temp[15] , \Add_add_temp[14] , \Add_add_temp[13] , 
            \Add_add_temp[12] , \Add_add_temp[11] , \Add_add_temp[10] , 
            \Add_add_temp[9] , \Add_add_temp[8] , \Add_add_temp[7] , \Add_add_temp[6] , 
            \Add_add_temp[5] , \Add_add_temp[4] , \Error_sub_temp[30] , 
            n19765, n14355, \qCurrent[3] , \qCurrent[4] , \qCurrent[5] , 
            \qCurrent[6] , \qCurrent[7] , \qCurrent[8] , \qCurrent[9] , 
            \qCurrent[10] , \qCurrent[11] , \qCurrent[12] , \qCurrent[13] , 
            \qCurrent[14] , \qCurrent[15] , \qCurrent[16] , \qCurrent[17] , 
            \qCurrent[18] , \qCurrent[19] , \qCurrent[20] , \qCurrent[21] , 
            \qCurrent[22] , \qCurrent[23] , \qCurrent[24] , \qCurrent[25] , 
            \qCurrent[26] , \qCurrent[27] , \qCurrent[28] , \qCurrent[29] , 
            \qCurrent[30] , \qCurrent[31] , n142, Saturate_out1_31__N_267, 
            Saturate_out1_31__N_266, Look_Up_Table_out1_1, n579, n17, 
            n267, n120, n14, n414, n11, n19604, n789, n785, 
            n781, n8, n777, n19351, n773, n769, n765, n270, 
            n123, n761, n757, n417, n753, n749, n745, n741, 
            n737, n489, n489_adj_32, n342, n342_adj_33, n246, n288, 
            n285, n282, n279, n276, n273, n258, n255, n252, 
            n261, n249, n44, n126, n420, n129, n423, n41, n86, 
            n89, n86_adj_34, n83, n80, n19702, n77, n74, n38, 
            n71, n68, n65, n62, n59, n56, n50, n53, n92, n244, 
            n35, n195, n114, n108, n102, n99, \Product2_mul_temp[2] , 
            n141_adj_35, n105, n138, n135, n132, n111, n32, n538, 
            n29, n426, n685, n402, n429, n432, n26, n391, n23, 
            n391_adj_36, n576, n576_adj_37, n573, n570, n567, n564, 
            n405, n628, n625, n622, n435, n619, n616, n613, 
            n610, n607, n601, n561, n598, n595, n592, n589, 
            n604, n631, n558, n20, n264, n117, n411, n587, n587_adj_38, 
            n582, n393, n408, n555, n552, n549, n396, n399, 
            n546, n543, n540, \Error_sub_temp[31]_adj_39 , n146_adj_40, 
            \preSatVoltage[23]_adj_41 , \preSatVoltage[19]_adj_42 , n794_adj_43, 
            \preSatVoltage[12]_adj_44 , n141_adj_45, \Error_sub_temp[30]_adj_46 , 
            Out_31__N_333_adj_47, Out_31__N_332_adj_48, \dVoltage[5] , 
            \dVoltage[2] , \dVoltage[8] , \dVoltage[12] , \dVoltage[15] , 
            \dVoltage[13] , \dVoltage[6] , \dVoltage[9] , \dVoltage[11] , 
            \dVoltage[10] , \dVoltage[7] , \dVoltage[3] , \dVoltage[14] , 
            \preSatVoltage[10]_adj_49 , n142_adj_50, n14349, n14348, 
            n14347, n14346, n14345, n14344, n14343, n14342, n14341, 
            n14340, n14339, n14338, n14320, n14337, n14336, n14335, 
            n14334, n14333, n14332, n14331, n14330, n14329, \Add_add_temp[34]_adj_51 , 
            \Add_add_temp[33]_adj_52 , \Add_add_temp[32]_adj_53 , \Add_add_temp[31]_adj_54 , 
            \Add_add_temp[30]_adj_55 , \Add_add_temp[29]_adj_56 , \Add_add_temp[28]_adj_57 , 
            \Add_add_temp[27]_adj_58 , \Add_add_temp[26]_adj_59 , \Add_add_temp[25]_adj_60 , 
            \Add_add_temp[24]_adj_61 , \Add_add_temp[23]_adj_62 , \Add_add_temp[22]_adj_63 , 
            \Add_add_temp[21]_adj_64 , \Add_add_temp[20]_adj_65 , \Add_add_temp[19]_adj_66 , 
            \Add_add_temp[18]_adj_67 , \Add_add_temp[17]_adj_68 , \Add_add_temp[16]_adj_69 , 
            \Add_add_temp[15]_adj_70 , \Add_add_temp[14]_adj_71 , \Add_add_temp[13]_adj_72 , 
            \Add_add_temp[12]_adj_73 , \Add_add_temp[11]_adj_74 , \Add_add_temp[10]_adj_75 , 
            \Add_add_temp[9]_adj_76 , \Add_add_temp[8]_adj_77 , \Add_add_temp[7]_adj_78 , 
            \Add_add_temp[6]_adj_79 , \Add_add_temp[5]_adj_80 , \Add_add_temp[4]_adj_81 , 
            n14328, n14327, n14326, n14322, n793_adj_82, n14325, 
            n19782, n14324, n14323, n14321, Saturate_out1_31__N_267_adj_83, 
            Saturate_out1_31__N_266_adj_84, \dCurrent[3] , \dCurrent[4] , 
            \dCurrent[5] , \dCurrent[6] , \dCurrent[7] , \dCurrent[8] , 
            \dCurrent[9] , \dCurrent[10] , \dCurrent[11] , \dCurrent[12] , 
            \dCurrent[13] , \dCurrent[14] , \dCurrent[15] , \dCurrent[16] , 
            \dCurrent[17] , \dCurrent[18] , \dCurrent[19] , \dCurrent[20] , 
            \dCurrent[21] , \dCurrent[22] , \dCurrent[23] , \dCurrent[24] , 
            \dCurrent[25] , \dCurrent[26] , \dCurrent[27] , \dCurrent[28] , 
            \dCurrent[29] , \dCurrent[30] , \dCurrent[31] , n342_adj_85, 
            n342_adj_86, n114_adj_87, n408_adj_88, n14_adj_89, n604_adj_90, 
            n685_adj_91, n685_adj_92, n417_adj_93, n123_adj_94, n613_adj_95, 
            n429_adj_96, n135_adj_97, n625_adj_98, n587_adj_99, n587_adj_100, 
            n399_adj_101, n426_adj_102, n414_adj_103, n432_adj_104, 
            n393_adj_105, n405_adj_106, n402_adj_107, n396_adj_108, 
            n420_adj_109, n423_adj_110, n44_adj_111, n489_adj_112, n8_adj_113, 
            n489_adj_114, n20_adj_115, n126_adj_116, n616_adj_117, n391_adj_118, 
            n391_adj_119, n19576, n129_adj_120, n619_adj_121, n11_adj_122, 
            n35_adj_123, n19352, n26_adj_124, \Product3_mul_temp[2] , 
            n120_adj_125, n111_adj_126, n102_adj_127, n99_adj_128, n108_adj_129, 
            n138_adj_130, n132_adj_131, n105_adj_132, n610_adj_133, 
            n595_adj_134, n23_adj_135, n622_adj_136, n41_adj_137, n601_adj_138, 
            n592_adj_139, n598_adj_140, n589_adj_141, n628_adj_142, 
            n32_adj_143, n538_adj_144, n29_adj_145, n17_adj_146, n71_adj_147, 
            n83_adj_148, n59_adj_149, n50_adj_150, n92_adj_151, n68_adj_152, 
            n62_adj_153, n53_adj_154, n65_adj_155, n38_adj_156, n56_adj_157, 
            n80_adj_158, n244_adj_159, n233, n200, n203, n86_adj_160, 
            n77_adj_161, n197, n239, n206, n86_adj_162, n215, n89_adj_163, 
            n74_adj_164, n227, n233_adj_165, n224, n221, n209, n236, 
            n230, n244_adj_166, n212, n218, n279_adj_167, n270_adj_168, 
            n267_adj_169, n255_adj_170, n285_adj_171, n264_adj_172, 
            n258_adj_173, n249_adj_174, n246_adj_175, n273_adj_176, 
            n282_adj_177, n261_adj_178, n19681, n288_adj_179, n276_adj_180, 
            n252_adj_181, n789_adj_182, n785_adj_183, n765_adj_184, 
            n753_adj_185, n741_adj_186, n757_adj_187, n745_adj_188, 
            n761_adj_189, n195_adj_190, n737_adj_191, n749_adj_192, 
            n781_adj_193, n777_adj_194, n773_adj_195, n769_adj_196, 
            n19684, n435_adj_197, n141_adj_198, n631_adj_199, n117_adj_200, 
            n411_adj_201, n607_adj_202) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n14381;
    input pin3_clk_16mhz_N_keep;
    input \Product_mul_temp[26] ;
    output \Error_sub_temp[31] ;
    output \preSatVoltage[10] ;
    output Out_31__N_333;
    output Out_31__N_332;
    output \qVoltage[8] ;
    output \qVoltage[5] ;
    output \qVoltage[2] ;
    output \qVoltage[12] ;
    input n14380;
    output \preSatVoltage[23] ;
    output \qVoltage[14] ;
    output \qVoltage[9] ;
    input n14379;
    output \preSatVoltage[13] ;
    output \preSatVoltage[12] ;
    output \qVoltage[4] ;
    output \qVoltage[3] ;
    output \qVoltage[15] ;
    input n14378;
    input n14377;
    input n14376;
    input n14375;
    input n14374;
    output \qVoltage[6] ;
    input n14373;
    output \preSatVoltage[22] ;
    output \preSatVoltage[19] ;
    output \qVoltage[13] ;
    output \qVoltage[10] ;
    output \qVoltage[7] ;
    input n14354;
    input n14372;
    input n14371;
    input n14370;
    input n14369;
    input n14353;
    input n14368;
    input n14367;
    input n14366;
    input n14365;
    input n14364;
    input n14363;
    input n14362;
    input n14361;
    input n14360;
    input n14359;
    input n14352;
    input n14358;
    input \Amp25_out1[14] ;
    output n146;
    input n14357;
    input n14356;
    input n793;
    input n141;
    input n794;
    output \Add_add_temp[34] ;
    output \Add_add_temp[33] ;
    output \Add_add_temp[32] ;
    output \Add_add_temp[31] ;
    output \Add_add_temp[30] ;
    output \Add_add_temp[29] ;
    output \Add_add_temp[28] ;
    output \Add_add_temp[27] ;
    output \Add_add_temp[26] ;
    output \Add_add_temp[25] ;
    output \Add_add_temp[24] ;
    output \Add_add_temp[23] ;
    output \Add_add_temp[22] ;
    output \Add_add_temp[21] ;
    output \Add_add_temp[20] ;
    output \Add_add_temp[19] ;
    output \Add_add_temp[18] ;
    output \Add_add_temp[17] ;
    output \Add_add_temp[16] ;
    output \Add_add_temp[15] ;
    output \Add_add_temp[14] ;
    output \Add_add_temp[13] ;
    output \Add_add_temp[12] ;
    output \Add_add_temp[11] ;
    output \Add_add_temp[10] ;
    output \Add_add_temp[9] ;
    output \Add_add_temp[8] ;
    output \Add_add_temp[7] ;
    output \Add_add_temp[6] ;
    output \Add_add_temp[5] ;
    output \Add_add_temp[4] ;
    output \Error_sub_temp[30] ;
    input n19765;
    input n14355;
    input \qCurrent[3] ;
    input \qCurrent[4] ;
    input \qCurrent[5] ;
    input \qCurrent[6] ;
    input \qCurrent[7] ;
    input \qCurrent[8] ;
    input \qCurrent[9] ;
    input \qCurrent[10] ;
    input \qCurrent[11] ;
    input \qCurrent[12] ;
    input \qCurrent[13] ;
    input \qCurrent[14] ;
    input \qCurrent[15] ;
    input \qCurrent[16] ;
    input \qCurrent[17] ;
    input \qCurrent[18] ;
    input \qCurrent[19] ;
    input \qCurrent[20] ;
    input \qCurrent[21] ;
    input \qCurrent[22] ;
    input \qCurrent[23] ;
    input \qCurrent[24] ;
    input \qCurrent[25] ;
    input \qCurrent[26] ;
    input \qCurrent[27] ;
    input \qCurrent[28] ;
    input \qCurrent[29] ;
    input \qCurrent[30] ;
    input \qCurrent[31] ;
    input n142;
    output Saturate_out1_31__N_267;
    output Saturate_out1_31__N_266;
    input [15:0]Look_Up_Table_out1_1;
    output n579;
    output n17;
    output n267;
    output n120;
    output n14;
    output n414;
    output n11;
    output n19604;
    output n789;
    output n785;
    output n781;
    output n8;
    output n777;
    output n19351;
    output n773;
    output n769;
    output n765;
    output n270;
    output n123;
    output n761;
    output n757;
    output n417;
    output n753;
    output n749;
    output n745;
    output n741;
    output n737;
    output n489;
    output n489_adj_32;
    output n342;
    output n342_adj_33;
    output n246;
    output n288;
    output n285;
    output n282;
    output n279;
    output n276;
    output n273;
    output n258;
    output n255;
    output n252;
    output n261;
    output n249;
    output n44;
    output n126;
    output n420;
    output n129;
    output n423;
    output n41;
    output n86;
    output n89;
    output n86_adj_34;
    output n83;
    output n80;
    output n19702;
    output n77;
    output n74;
    output n38;
    output n71;
    output n68;
    output n65;
    output n62;
    output n59;
    output n56;
    output n50;
    output n53;
    output n92;
    output n244;
    output n35;
    output n195;
    output n114;
    output n108;
    output n102;
    output n99;
    output \Product2_mul_temp[2] ;
    output n141_adj_35;
    output n105;
    output n138;
    output n135;
    output n132;
    output n111;
    output n32;
    output n538;
    output n29;
    output n426;
    output n685;
    output n402;
    output n429;
    output n432;
    output n26;
    output n391;
    output n23;
    output n391_adj_36;
    output n576;
    output n576_adj_37;
    output n573;
    output n570;
    output n567;
    output n564;
    output n405;
    output n628;
    output n625;
    output n622;
    output n435;
    output n619;
    output n616;
    output n613;
    output n610;
    output n607;
    output n601;
    output n561;
    output n598;
    output n595;
    output n592;
    output n589;
    output n604;
    output n631;
    output n558;
    output n20;
    output n264;
    output n117;
    output n411;
    output n587;
    output n587_adj_38;
    output n582;
    output n393;
    output n408;
    output n555;
    output n552;
    output n549;
    output n396;
    output n399;
    output n546;
    output n543;
    output n540;
    output \Error_sub_temp[31]_adj_39 ;
    output n146_adj_40;
    output \preSatVoltage[23]_adj_41 ;
    output \preSatVoltage[19]_adj_42 ;
    input n794_adj_43;
    output \preSatVoltage[12]_adj_44 ;
    input n141_adj_45;
    output \Error_sub_temp[30]_adj_46 ;
    output Out_31__N_333_adj_47;
    output Out_31__N_332_adj_48;
    output \dVoltage[5] ;
    output \dVoltage[2] ;
    output \dVoltage[8] ;
    output \dVoltage[12] ;
    output \dVoltage[15] ;
    output \dVoltage[13] ;
    output \dVoltage[6] ;
    output \dVoltage[9] ;
    output \dVoltage[11] ;
    output \dVoltage[10] ;
    output \dVoltage[7] ;
    output \dVoltage[3] ;
    output \dVoltage[14] ;
    output \preSatVoltage[10]_adj_49 ;
    input n142_adj_50;
    input n14349;
    input n14348;
    input n14347;
    input n14346;
    input n14345;
    input n14344;
    input n14343;
    input n14342;
    input n14341;
    input n14340;
    input n14339;
    input n14338;
    input n14320;
    input n14337;
    input n14336;
    input n14335;
    input n14334;
    input n14333;
    input n14332;
    input n14331;
    input n14330;
    input n14329;
    output \Add_add_temp[34]_adj_51 ;
    output \Add_add_temp[33]_adj_52 ;
    output \Add_add_temp[32]_adj_53 ;
    output \Add_add_temp[31]_adj_54 ;
    output \Add_add_temp[30]_adj_55 ;
    output \Add_add_temp[29]_adj_56 ;
    output \Add_add_temp[28]_adj_57 ;
    output \Add_add_temp[27]_adj_58 ;
    output \Add_add_temp[26]_adj_59 ;
    output \Add_add_temp[25]_adj_60 ;
    output \Add_add_temp[24]_adj_61 ;
    output \Add_add_temp[23]_adj_62 ;
    output \Add_add_temp[22]_adj_63 ;
    output \Add_add_temp[21]_adj_64 ;
    output \Add_add_temp[20]_adj_65 ;
    output \Add_add_temp[19]_adj_66 ;
    output \Add_add_temp[18]_adj_67 ;
    output \Add_add_temp[17]_adj_68 ;
    output \Add_add_temp[16]_adj_69 ;
    output \Add_add_temp[15]_adj_70 ;
    output \Add_add_temp[14]_adj_71 ;
    output \Add_add_temp[13]_adj_72 ;
    output \Add_add_temp[12]_adj_73 ;
    output \Add_add_temp[11]_adj_74 ;
    output \Add_add_temp[10]_adj_75 ;
    output \Add_add_temp[9]_adj_76 ;
    output \Add_add_temp[8]_adj_77 ;
    output \Add_add_temp[7]_adj_78 ;
    output \Add_add_temp[6]_adj_79 ;
    output \Add_add_temp[5]_adj_80 ;
    output \Add_add_temp[4]_adj_81 ;
    input n14328;
    input n14327;
    input n14326;
    input n14322;
    input n793_adj_82;
    input n14325;
    input n19782;
    input n14324;
    input n14323;
    input n14321;
    output Saturate_out1_31__N_267_adj_83;
    output Saturate_out1_31__N_266_adj_84;
    input \dCurrent[3] ;
    input \dCurrent[4] ;
    input \dCurrent[5] ;
    input \dCurrent[6] ;
    input \dCurrent[7] ;
    input \dCurrent[8] ;
    input \dCurrent[9] ;
    input \dCurrent[10] ;
    input \dCurrent[11] ;
    input \dCurrent[12] ;
    input \dCurrent[13] ;
    input \dCurrent[14] ;
    input \dCurrent[15] ;
    input \dCurrent[16] ;
    input \dCurrent[17] ;
    input \dCurrent[18] ;
    input \dCurrent[19] ;
    input \dCurrent[20] ;
    input \dCurrent[21] ;
    input \dCurrent[22] ;
    input \dCurrent[23] ;
    input \dCurrent[24] ;
    input \dCurrent[25] ;
    input \dCurrent[26] ;
    input \dCurrent[27] ;
    input \dCurrent[28] ;
    input \dCurrent[29] ;
    input \dCurrent[30] ;
    input \dCurrent[31] ;
    output n342_adj_85;
    output n342_adj_86;
    output n114_adj_87;
    output n408_adj_88;
    output n14_adj_89;
    output n604_adj_90;
    output n685_adj_91;
    output n685_adj_92;
    output n417_adj_93;
    output n123_adj_94;
    output n613_adj_95;
    output n429_adj_96;
    output n135_adj_97;
    output n625_adj_98;
    output n587_adj_99;
    output n587_adj_100;
    output n399_adj_101;
    output n426_adj_102;
    output n414_adj_103;
    output n432_adj_104;
    output n393_adj_105;
    output n405_adj_106;
    output n402_adj_107;
    output n396_adj_108;
    output n420_adj_109;
    output n423_adj_110;
    output n44_adj_111;
    output n489_adj_112;
    output n8_adj_113;
    output n489_adj_114;
    output n20_adj_115;
    output n126_adj_116;
    output n616_adj_117;
    output n391_adj_118;
    output n391_adj_119;
    output n19576;
    output n129_adj_120;
    output n619_adj_121;
    output n11_adj_122;
    output n35_adj_123;
    output n19352;
    output n26_adj_124;
    output \Product3_mul_temp[2] ;
    output n120_adj_125;
    output n111_adj_126;
    output n102_adj_127;
    output n99_adj_128;
    output n108_adj_129;
    output n138_adj_130;
    output n132_adj_131;
    output n105_adj_132;
    output n610_adj_133;
    output n595_adj_134;
    output n23_adj_135;
    output n622_adj_136;
    output n41_adj_137;
    output n601_adj_138;
    output n592_adj_139;
    output n598_adj_140;
    output n589_adj_141;
    output n628_adj_142;
    output n32_adj_143;
    output n538_adj_144;
    output n29_adj_145;
    output n17_adj_146;
    output n71_adj_147;
    output n83_adj_148;
    output n59_adj_149;
    output n50_adj_150;
    output n92_adj_151;
    output n68_adj_152;
    output n62_adj_153;
    output n53_adj_154;
    output n65_adj_155;
    output n38_adj_156;
    output n56_adj_157;
    output n80_adj_158;
    output n244_adj_159;
    output n233;
    output n200;
    output n203;
    output n86_adj_160;
    output n77_adj_161;
    output n197;
    output n239;
    output n206;
    output n86_adj_162;
    output n215;
    output n89_adj_163;
    output n74_adj_164;
    output n227;
    output n233_adj_165;
    output n224;
    output n221;
    output n209;
    output n236;
    output n230;
    output n244_adj_166;
    output n212;
    output n218;
    output n279_adj_167;
    output n270_adj_168;
    output n267_adj_169;
    output n255_adj_170;
    output n285_adj_171;
    output n264_adj_172;
    output n258_adj_173;
    output n249_adj_174;
    output n246_adj_175;
    output n273_adj_176;
    output n282_adj_177;
    output n261_adj_178;
    output n19681;
    output n288_adj_179;
    output n276_adj_180;
    output n252_adj_181;
    output n789_adj_182;
    output n785_adj_183;
    output n765_adj_184;
    output n753_adj_185;
    output n741_adj_186;
    output n757_adj_187;
    output n745_adj_188;
    output n761_adj_189;
    output n195_adj_190;
    output n737_adj_191;
    output n749_adj_192;
    output n781_adj_193;
    output n777_adj_194;
    output n773_adj_195;
    output n769_adj_196;
    output n19684;
    output n435_adj_197;
    output n141_adj_198;
    output n631_adj_199;
    output n117_adj_200;
    output n411_adj_201;
    output n607_adj_202;
    
    wire [29:0]n1;
    
    D_Current_Control u_Q_Current_Control (.GND_net(GND_net), .n14381(n14381), 
            .pin3_clk_16mhz_N_keep(pin3_clk_16mhz_N_keep), .\Product_mul_temp[26] (\Product_mul_temp[26] ), 
            .\Error_sub_temp[31] (\Error_sub_temp[31] ), .\preSatVoltage[10] (\preSatVoltage[10] ), 
            .Out_31__N_333(Out_31__N_333), .Out_31__N_332(Out_31__N_332), 
            .\qVoltage[8] (\qVoltage[8] ), .\qVoltage[5] (\qVoltage[5] ), 
            .\qVoltage[2] (\qVoltage[2] ), .\qVoltage[12] (\qVoltage[12] ), 
            .n14380(n14380), .\preSatVoltage[23] (\preSatVoltage[23] ), 
            .\qVoltage[14] (\qVoltage[14] ), .\qVoltage[9] (\qVoltage[9] ), 
            .n14379(n14379), .\preSatVoltage[13] (\preSatVoltage[13] ), 
            .\preSatVoltage[12] (\preSatVoltage[12] ), .\qVoltage[4] (\qVoltage[4] ), 
            .\qVoltage[3] (\qVoltage[3] ), .\qVoltage[15] (\qVoltage[15] ), 
            .n14378(n14378), .n14377(n14377), .n14376(n14376), .n14375(n14375), 
            .n14374(n14374), .\qVoltage[6] (\qVoltage[6] ), .n14373(n14373), 
            .\preSatVoltage[22] (\preSatVoltage[22] ), .\preSatVoltage[19] (\preSatVoltage[19] ), 
            .\qVoltage[13] (\qVoltage[13] ), .\qVoltage[10] (\qVoltage[10] ), 
            .\qVoltage[7] (\qVoltage[7] ), .n14354(n14354), .n14372(n14372), 
            .n14371(n14371), .n14370(n14370), .n14369(n14369), .n14353(n14353), 
            .n14368(n14368), .n14367(n14367), .n14366(n14366), .n14365(n14365), 
            .n14364(n14364), .n14363(n14363), .n14362(n14362), .n14361(n14361), 
            .n14360(n14360), .n14359(n14359), .n14352(n14352), .n14358(n14358), 
            .\Amp25_out1[14] (\Amp25_out1[14] ), .n146(n146), .n14357(n14357), 
            .n14356(n14356), .n793(n793), .n141(n141), .n794(n794), 
            .\Add_add_temp[34] (\Add_add_temp[34] ), .\Add_add_temp[33] (\Add_add_temp[33] ), 
            .\Add_add_temp[32] (\Add_add_temp[32] ), .\Add_add_temp[31] (\Add_add_temp[31] ), 
            .\Add_add_temp[30] (\Add_add_temp[30] ), .\Add_add_temp[29] (\Add_add_temp[29] ), 
            .\Add_add_temp[28] (\Add_add_temp[28] ), .\Add_add_temp[27] (\Add_add_temp[27] ), 
            .\Add_add_temp[26] (\Add_add_temp[26] ), .\Add_add_temp[25] (\Add_add_temp[25] ), 
            .\Add_add_temp[24] (\Add_add_temp[24] ), .\Add_add_temp[23] (\Add_add_temp[23] ), 
            .\Add_add_temp[22] (\Add_add_temp[22] ), .\Add_add_temp[21] (\Add_add_temp[21] ), 
            .\Add_add_temp[20] (\Add_add_temp[20] ), .\Add_add_temp[19] (\Add_add_temp[19] ), 
            .\Add_add_temp[18] (\Add_add_temp[18] ), .\Add_add_temp[17] (\Add_add_temp[17] ), 
            .\Add_add_temp[16] (\Add_add_temp[16] ), .\Add_add_temp[15] (\Add_add_temp[15] ), 
            .\Add_add_temp[14] (\Add_add_temp[14] ), .\Add_add_temp[13] (\Add_add_temp[13] ), 
            .\Add_add_temp[12] (\Add_add_temp[12] ), .\Add_add_temp[11] (\Add_add_temp[11] ), 
            .\Add_add_temp[10] (\Add_add_temp[10] ), .\Add_add_temp[9] (\Add_add_temp[9] ), 
            .\Add_add_temp[8] (\Add_add_temp[8] ), .\Add_add_temp[7] (\Add_add_temp[7] ), 
            .\Add_add_temp[6] (\Add_add_temp[6] ), .\Add_add_temp[5] (\Add_add_temp[5] ), 
            .\Add_add_temp[4] (\Add_add_temp[4] ), .\Error_sub_temp[30] (\Error_sub_temp[30] ), 
            .n31(n1[0]), .n19765(n19765), .n14355(n14355), .\qCurrent[3] (\qCurrent[3] ), 
            .\qCurrent[4] (\qCurrent[4] ), .\qCurrent[5] (\qCurrent[5] ), 
            .\qCurrent[6] (\qCurrent[6] ), .\qCurrent[7] (\qCurrent[7] ), 
            .\qCurrent[8] (\qCurrent[8] ), .\qCurrent[9] (\qCurrent[9] ), 
            .\qCurrent[10] (\qCurrent[10] ), .\qCurrent[11] (\qCurrent[11] ), 
            .\qCurrent[12] (\qCurrent[12] ), .\qCurrent[13] (\qCurrent[13] ), 
            .\qCurrent[14] (\qCurrent[14] ), .\qCurrent[15] (\qCurrent[15] ), 
            .\qCurrent[16] (\qCurrent[16] ), .\qCurrent[17] (\qCurrent[17] ), 
            .\qCurrent[18] (\qCurrent[18] ), .\qCurrent[19] (\qCurrent[19] ), 
            .\qCurrent[20] (\qCurrent[20] ), .\qCurrent[21] (\qCurrent[21] ), 
            .\qCurrent[22] (\qCurrent[22] ), .\qCurrent[23] (\qCurrent[23] ), 
            .\qCurrent[24] (\qCurrent[24] ), .\qCurrent[25] (\qCurrent[25] ), 
            .\qCurrent[26] (\qCurrent[26] ), .\qCurrent[27] (\qCurrent[27] ), 
            .\qCurrent[28] (\qCurrent[28] ), .\qCurrent[29] (\qCurrent[29] ), 
            .\qCurrent[30] (\qCurrent[30] ), .\qCurrent[31] (\qCurrent[31] ), 
            .n142(n142), .Saturate_out1_31__N_267(Saturate_out1_31__N_267), 
            .Saturate_out1_31__N_266(Saturate_out1_31__N_266), .Look_Up_Table_out1_1({Look_Up_Table_out1_1}), 
            .n579(n579), .n17(n17), .n267(n267), .n120(n120), .n14(n14), 
            .n414(n414), .n11(n11), .n19604(n19604), .n789(n789), .n785(n785), 
            .n781(n781), .n8(n8), .n777(n777), .n19351(n19351), .n773(n773), 
            .n769(n769), .n765(n765), .n270(n270), .n123(n123), .n761(n761), 
            .n757(n757), .n417(n417), .n753(n753), .n749(n749), .n745(n745), 
            .n741(n741), .n737(n737), .n489(n489), .n489_adj_25(n489_adj_32), 
            .n342(n342), .n342_adj_26(n342_adj_33), .n246(n246), .n288(n288), 
            .n285(n285), .n282(n282), .n279(n279), .n276(n276), .n273(n273), 
            .n258(n258), .n255(n255), .n252(n252), .n261(n261), .n249(n249), 
            .n44(n44), .n126(n126), .n420(n420), .n129(n129), .n423(n423), 
            .n41(n41), .n86(n86), .n89(n89), .n86_adj_27(n86_adj_34), 
            .n83(n83), .n80(n80), .n19702(n19702), .n77(n77), .n74(n74), 
            .n38(n38), .n71(n71), .n68(n68), .n65(n65), .n62(n62), 
            .n59(n59), .n56(n56), .n50(n50), .n53(n53), .n92(n92), 
            .n244(n244), .n35(n35), .n195(n195), .n114(n114), .n108(n108), 
            .n102(n102), .n99(n99), .\Product2_mul_temp[2] (\Product2_mul_temp[2] ), 
            .n141_adj_28(n141_adj_35), .n105(n105), .n138(n138), .n135(n135), 
            .n132(n132), .n111(n111), .n32(n32), .n538(n538), .n29(n29), 
            .n426(n426), .n685(n685), .n402(n402), .n429(n429), .n432(n432), 
            .n26(n26), .n391(n391), .n23(n23), .n391_adj_29(n391_adj_36), 
            .n576(n576), .n576_adj_30(n576_adj_37), .n573(n573), .n570(n570), 
            .n567(n567), .n564(n564), .n405(n405), .n628(n628), .n625(n625), 
            .n622(n622), .n435(n435), .n619(n619), .n616(n616), .n613(n613), 
            .n610(n610), .n607(n607), .n601(n601), .n561(n561), .n598(n598), 
            .n595(n595), .n592(n592), .n589(n589), .n604(n604), .n631(n631), 
            .n558(n558), .n20(n20), .n264(n264), .n117(n117), .n411(n411), 
            .n587(n587), .n587_adj_31(n587_adj_38), .n582(n582), .n393(n393), 
            .n408(n408), .n555(n555), .n552(n552), .n549(n549), .n396(n396), 
            .n399(n399), .n546(n546), .n543(n543), .n540(n540)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/DQ_Current_Control.v(67[21] 75[43])
    D_Current_Control_U1 u_D_Current_Control (.GND_net(GND_net), .\Product_mul_temp[26] (\Product_mul_temp[26] ), 
            .\Error_sub_temp[31] (\Error_sub_temp[31]_adj_39 ), .n146(n146_adj_40), 
            .\preSatVoltage[23] (\preSatVoltage[23]_adj_41 ), .\preSatVoltage[19] (\preSatVoltage[19]_adj_42 ), 
            .n794(n794_adj_43), .pin3_clk_16mhz_N_keep(pin3_clk_16mhz_N_keep), 
            .\preSatVoltage[12] (\preSatVoltage[12]_adj_44 ), .n141(n141_adj_45), 
            .\Error_sub_temp[30] (\Error_sub_temp[30]_adj_46 ), .Out_31__N_333(Out_31__N_333_adj_47), 
            .Out_31__N_332(Out_31__N_332_adj_48), .\dVoltage[5] (\dVoltage[5] ), 
            .\dVoltage[2] (\dVoltage[2] ), .\dVoltage[8] (\dVoltage[8] ), 
            .\dVoltage[12] (\dVoltage[12] ), .\dVoltage[15] (\dVoltage[15] ), 
            .\dVoltage[13] (\dVoltage[13] ), .\dVoltage[6] (\dVoltage[6] ), 
            .\dVoltage[9] (\dVoltage[9] ), .\dVoltage[11] (\dVoltage[11] ), 
            .\dVoltage[10] (\dVoltage[10] ), .\dVoltage[7] (\dVoltage[7] ), 
            .\dVoltage[3] (\dVoltage[3] ), .\dVoltage[14] (\dVoltage[14] ), 
            .\preSatVoltage[10] (\preSatVoltage[10]_adj_49 ), .n142(n142_adj_50), 
            .n14349(n14349), .n14348(n14348), .n14347(n14347), .n14346(n14346), 
            .n14345(n14345), .n14344(n14344), .n14343(n14343), .n14342(n14342), 
            .n14341(n14341), .n14340(n14340), .n14339(n14339), .n14338(n14338), 
            .n14320(n14320), .n14337(n14337), .n14336(n14336), .n14335(n14335), 
            .n14334(n14334), .n14333(n14333), .n14332(n14332), .n14331(n14331), 
            .n14330(n14330), .n14329(n14329), .\Add_add_temp[34] (\Add_add_temp[34]_adj_51 ), 
            .\Add_add_temp[33] (\Add_add_temp[33]_adj_52 ), .\Add_add_temp[32] (\Add_add_temp[32]_adj_53 ), 
            .\Add_add_temp[31] (\Add_add_temp[31]_adj_54 ), .\Add_add_temp[30] (\Add_add_temp[30]_adj_55 ), 
            .\Add_add_temp[29] (\Add_add_temp[29]_adj_56 ), .\Add_add_temp[28] (\Add_add_temp[28]_adj_57 ), 
            .\Add_add_temp[27] (\Add_add_temp[27]_adj_58 ), .\Add_add_temp[26] (\Add_add_temp[26]_adj_59 ), 
            .\Add_add_temp[25] (\Add_add_temp[25]_adj_60 ), .\Add_add_temp[24] (\Add_add_temp[24]_adj_61 ), 
            .\Add_add_temp[23] (\Add_add_temp[23]_adj_62 ), .\Add_add_temp[22] (\Add_add_temp[22]_adj_63 ), 
            .\Add_add_temp[21] (\Add_add_temp[21]_adj_64 ), .\Add_add_temp[20] (\Add_add_temp[20]_adj_65 ), 
            .\Add_add_temp[19] (\Add_add_temp[19]_adj_66 ), .\Add_add_temp[18] (\Add_add_temp[18]_adj_67 ), 
            .\Add_add_temp[17] (\Add_add_temp[17]_adj_68 ), .\Add_add_temp[16] (\Add_add_temp[16]_adj_69 ), 
            .\Add_add_temp[15] (\Add_add_temp[15]_adj_70 ), .\Add_add_temp[14] (\Add_add_temp[14]_adj_71 ), 
            .\Add_add_temp[13] (\Add_add_temp[13]_adj_72 ), .\Add_add_temp[12] (\Add_add_temp[12]_adj_73 ), 
            .\Add_add_temp[11] (\Add_add_temp[11]_adj_74 ), .\Add_add_temp[10] (\Add_add_temp[10]_adj_75 ), 
            .\Add_add_temp[9] (\Add_add_temp[9]_adj_76 ), .\Add_add_temp[8] (\Add_add_temp[8]_adj_77 ), 
            .\Add_add_temp[7] (\Add_add_temp[7]_adj_78 ), .\Add_add_temp[6] (\Add_add_temp[6]_adj_79 ), 
            .\Add_add_temp[5] (\Add_add_temp[5]_adj_80 ), .\Add_add_temp[4] (\Add_add_temp[4]_adj_81 ), 
            .n14328(n14328), .n14327(n14327), .n14326(n14326), .n14322(n14322), 
            .n793(n793_adj_82), .n14325(n14325), .n19782(n19782), .n14324(n14324), 
            .n31(n1[0]), .n14323(n14323), .n14321(n14321), .Saturate_out1_31__N_267(Saturate_out1_31__N_267_adj_83), 
            .Saturate_out1_31__N_266(Saturate_out1_31__N_266_adj_84), .\dCurrent[3] (\dCurrent[3] ), 
            .\dCurrent[4] (\dCurrent[4] ), .\dCurrent[5] (\dCurrent[5] ), 
            .\dCurrent[6] (\dCurrent[6] ), .\dCurrent[7] (\dCurrent[7] ), 
            .\dCurrent[8] (\dCurrent[8] ), .\dCurrent[9] (\dCurrent[9] ), 
            .\dCurrent[10] (\dCurrent[10] ), .\dCurrent[11] (\dCurrent[11] ), 
            .\dCurrent[12] (\dCurrent[12] ), .\dCurrent[13] (\dCurrent[13] ), 
            .\dCurrent[14] (\dCurrent[14] ), .\dCurrent[15] (\dCurrent[15] ), 
            .\dCurrent[16] (\dCurrent[16] ), .\dCurrent[17] (\dCurrent[17] ), 
            .\dCurrent[18] (\dCurrent[18] ), .\dCurrent[19] (\dCurrent[19] ), 
            .\dCurrent[20] (\dCurrent[20] ), .\dCurrent[21] (\dCurrent[21] ), 
            .\dCurrent[22] (\dCurrent[22] ), .\dCurrent[23] (\dCurrent[23] ), 
            .\dCurrent[24] (\dCurrent[24] ), .\dCurrent[25] (\dCurrent[25] ), 
            .\dCurrent[26] (\dCurrent[26] ), .\dCurrent[27] (\dCurrent[27] ), 
            .\dCurrent[28] (\dCurrent[28] ), .\dCurrent[29] (\dCurrent[29] ), 
            .\dCurrent[30] (\dCurrent[30] ), .\dCurrent[31] (\dCurrent[31] ), 
            .n342(n342_adj_85), .Look_Up_Table_out1_1({Look_Up_Table_out1_1}), 
            .n342_adj_10(n342_adj_86), .n114(n114_adj_87), .n408(n408_adj_88), 
            .n14(n14_adj_89), .n604(n604_adj_90), .n685(n685_adj_91), 
            .n685_adj_11(n685_adj_92), .n417(n417_adj_93), .n123(n123_adj_94), 
            .n613(n613_adj_95), .n429(n429_adj_96), .n135(n135_adj_97), 
            .n625(n625_adj_98), .n587(n587_adj_99), .n587_adj_12(n587_adj_100), 
            .n399(n399_adj_101), .n426(n426_adj_102), .n414(n414_adj_103), 
            .n432(n432_adj_104), .n393(n393_adj_105), .n405(n405_adj_106), 
            .n402(n402_adj_107), .n396(n396_adj_108), .n420(n420_adj_109), 
            .n423(n423_adj_110), .n44(n44_adj_111), .n489(n489_adj_112), 
            .n8(n8_adj_113), .n489_adj_13(n489_adj_114), .n20(n20_adj_115), 
            .n126(n126_adj_116), .n616(n616_adj_117), .n391(n391_adj_118), 
            .n391_adj_14(n391_adj_119), .n19576(n19576), .n129(n129_adj_120), 
            .n619(n619_adj_121), .n11(n11_adj_122), .n35(n35_adj_123), 
            .n19352(n19352), .n26(n26_adj_124), .\Product3_mul_temp[2] (\Product3_mul_temp[2] ), 
            .n120(n120_adj_125), .n111(n111_adj_126), .n102(n102_adj_127), 
            .n99(n99_adj_128), .n108(n108_adj_129), .n138(n138_adj_130), 
            .n132(n132_adj_131), .n105(n105_adj_132), .n610(n610_adj_133), 
            .n595(n595_adj_134), .n23(n23_adj_135), .n622(n622_adj_136), 
            .n41(n41_adj_137), .n601(n601_adj_138), .n592(n592_adj_139), 
            .n598(n598_adj_140), .n589(n589_adj_141), .n628(n628_adj_142), 
            .n32(n32_adj_143), .n538(n538_adj_144), .n29(n29_adj_145), 
            .n17(n17_adj_146), .n71(n71_adj_147), .n83(n83_adj_148), .n59(n59_adj_149), 
            .n50(n50_adj_150), .n92(n92_adj_151), .n68(n68_adj_152), .n62(n62_adj_153), 
            .n53(n53_adj_154), .n65(n65_adj_155), .n38(n38_adj_156), .n56(n56_adj_157), 
            .n80(n80_adj_158), .n244(n244_adj_159), .n233(n233), .n200(n200), 
            .n203(n203), .n86(n86_adj_160), .n77(n77_adj_161), .n197(n197), 
            .n239(n239), .n206(n206), .n86_adj_15(n86_adj_162), .n215(n215), 
            .n89(n89_adj_163), .n74(n74_adj_164), .n227(n227), .n233_adj_16(n233_adj_165), 
            .n224(n224), .n221(n221), .n209(n209), .n236(n236), .n230(n230), 
            .n244_adj_17(n244_adj_166), .n212(n212), .n218(n218), .n279(n279_adj_167), 
            .n270(n270_adj_168), .n267(n267_adj_169), .n255(n255_adj_170), 
            .n285(n285_adj_171), .n264(n264_adj_172), .n258(n258_adj_173), 
            .n249(n249_adj_174), .n246(n246_adj_175), .n273(n273_adj_176), 
            .n282(n282_adj_177), .n261(n261_adj_178), .n19681(n19681), 
            .n288(n288_adj_179), .n276(n276_adj_180), .n252(n252_adj_181), 
            .n789(n789_adj_182), .n785(n785_adj_183), .n765(n765_adj_184), 
            .n753(n753_adj_185), .n741(n741_adj_186), .n757(n757_adj_187), 
            .n745(n745_adj_188), .n761(n761_adj_189), .n195(n195_adj_190), 
            .n737(n737_adj_191), .n749(n749_adj_192), .n781(n781_adj_193), 
            .n777(n777_adj_194), .n773(n773_adj_195), .n769(n769_adj_196), 
            .n19684(n19684), .n435(n435_adj_197), .n141_adj_18(n141_adj_198), 
            .n631(n631_adj_199), .n117(n117_adj_200), .n411(n411_adj_201), 
            .n607(n607_adj_202)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/DQ_Current_Control.v(55[21] 63[43])
    
endmodule
//
// Verilog Description of module D_Current_Control
//

module D_Current_Control (GND_net, n14381, pin3_clk_16mhz_N_keep, \Product_mul_temp[26] , 
            \Error_sub_temp[31] , \preSatVoltage[10] , Out_31__N_333, 
            Out_31__N_332, \qVoltage[8] , \qVoltage[5] , \qVoltage[2] , 
            \qVoltage[12] , n14380, \preSatVoltage[23] , \qVoltage[14] , 
            \qVoltage[9] , n14379, \preSatVoltage[13] , \preSatVoltage[12] , 
            \qVoltage[4] , \qVoltage[3] , \qVoltage[15] , n14378, n14377, 
            n14376, n14375, n14374, \qVoltage[6] , n14373, \preSatVoltage[22] , 
            \preSatVoltage[19] , \qVoltage[13] , \qVoltage[10] , \qVoltage[7] , 
            n14354, n14372, n14371, n14370, n14369, n14353, n14368, 
            n14367, n14366, n14365, n14364, n14363, n14362, n14361, 
            n14360, n14359, n14352, n14358, \Amp25_out1[14] , n146, 
            n14357, n14356, n793, n141, n794, \Add_add_temp[34] , 
            \Add_add_temp[33] , \Add_add_temp[32] , \Add_add_temp[31] , 
            \Add_add_temp[30] , \Add_add_temp[29] , \Add_add_temp[28] , 
            \Add_add_temp[27] , \Add_add_temp[26] , \Add_add_temp[25] , 
            \Add_add_temp[24] , \Add_add_temp[23] , \Add_add_temp[22] , 
            \Add_add_temp[21] , \Add_add_temp[20] , \Add_add_temp[19] , 
            \Add_add_temp[18] , \Add_add_temp[17] , \Add_add_temp[16] , 
            \Add_add_temp[15] , \Add_add_temp[14] , \Add_add_temp[13] , 
            \Add_add_temp[12] , \Add_add_temp[11] , \Add_add_temp[10] , 
            \Add_add_temp[9] , \Add_add_temp[8] , \Add_add_temp[7] , \Add_add_temp[6] , 
            \Add_add_temp[5] , \Add_add_temp[4] , \Error_sub_temp[30] , 
            n31, n19765, n14355, \qCurrent[3] , \qCurrent[4] , \qCurrent[5] , 
            \qCurrent[6] , \qCurrent[7] , \qCurrent[8] , \qCurrent[9] , 
            \qCurrent[10] , \qCurrent[11] , \qCurrent[12] , \qCurrent[13] , 
            \qCurrent[14] , \qCurrent[15] , \qCurrent[16] , \qCurrent[17] , 
            \qCurrent[18] , \qCurrent[19] , \qCurrent[20] , \qCurrent[21] , 
            \qCurrent[22] , \qCurrent[23] , \qCurrent[24] , \qCurrent[25] , 
            \qCurrent[26] , \qCurrent[27] , \qCurrent[28] , \qCurrent[29] , 
            \qCurrent[30] , \qCurrent[31] , n142, Saturate_out1_31__N_267, 
            Saturate_out1_31__N_266, Look_Up_Table_out1_1, n579, n17, 
            n267, n120, n14, n414, n11, n19604, n789, n785, 
            n781, n8, n777, n19351, n773, n769, n765, n270, 
            n123, n761, n757, n417, n753, n749, n745, n741, 
            n737, n489, n489_adj_25, n342, n342_adj_26, n246, n288, 
            n285, n282, n279, n276, n273, n258, n255, n252, 
            n261, n249, n44, n126, n420, n129, n423, n41, n86, 
            n89, n86_adj_27, n83, n80, n19702, n77, n74, n38, 
            n71, n68, n65, n62, n59, n56, n50, n53, n92, n244, 
            n35, n195, n114, n108, n102, n99, \Product2_mul_temp[2] , 
            n141_adj_28, n105, n138, n135, n132, n111, n32, n538, 
            n29, n426, n685, n402, n429, n432, n26, n391, n23, 
            n391_adj_29, n576, n576_adj_30, n573, n570, n567, n564, 
            n405, n628, n625, n622, n435, n619, n616, n613, 
            n610, n607, n601, n561, n598, n595, n592, n589, 
            n604, n631, n558, n20, n264, n117, n411, n587, n587_adj_31, 
            n582, n393, n408, n555, n552, n549, n396, n399, 
            n546, n543, n540) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n14381;
    input pin3_clk_16mhz_N_keep;
    input \Product_mul_temp[26] ;
    output \Error_sub_temp[31] ;
    output \preSatVoltage[10] ;
    output Out_31__N_333;
    output Out_31__N_332;
    output \qVoltage[8] ;
    output \qVoltage[5] ;
    output \qVoltage[2] ;
    output \qVoltage[12] ;
    input n14380;
    output \preSatVoltage[23] ;
    output \qVoltage[14] ;
    output \qVoltage[9] ;
    input n14379;
    output \preSatVoltage[13] ;
    output \preSatVoltage[12] ;
    output \qVoltage[4] ;
    output \qVoltage[3] ;
    output \qVoltage[15] ;
    input n14378;
    input n14377;
    input n14376;
    input n14375;
    input n14374;
    output \qVoltage[6] ;
    input n14373;
    output \preSatVoltage[22] ;
    output \preSatVoltage[19] ;
    output \qVoltage[13] ;
    output \qVoltage[10] ;
    output \qVoltage[7] ;
    input n14354;
    input n14372;
    input n14371;
    input n14370;
    input n14369;
    input n14353;
    input n14368;
    input n14367;
    input n14366;
    input n14365;
    input n14364;
    input n14363;
    input n14362;
    input n14361;
    input n14360;
    input n14359;
    input n14352;
    input n14358;
    input \Amp25_out1[14] ;
    output n146;
    input n14357;
    input n14356;
    input n793;
    input n141;
    input n794;
    output \Add_add_temp[34] ;
    output \Add_add_temp[33] ;
    output \Add_add_temp[32] ;
    output \Add_add_temp[31] ;
    output \Add_add_temp[30] ;
    output \Add_add_temp[29] ;
    output \Add_add_temp[28] ;
    output \Add_add_temp[27] ;
    output \Add_add_temp[26] ;
    output \Add_add_temp[25] ;
    output \Add_add_temp[24] ;
    output \Add_add_temp[23] ;
    output \Add_add_temp[22] ;
    output \Add_add_temp[21] ;
    output \Add_add_temp[20] ;
    output \Add_add_temp[19] ;
    output \Add_add_temp[18] ;
    output \Add_add_temp[17] ;
    output \Add_add_temp[16] ;
    output \Add_add_temp[15] ;
    output \Add_add_temp[14] ;
    output \Add_add_temp[13] ;
    output \Add_add_temp[12] ;
    output \Add_add_temp[11] ;
    output \Add_add_temp[10] ;
    output \Add_add_temp[9] ;
    output \Add_add_temp[8] ;
    output \Add_add_temp[7] ;
    output \Add_add_temp[6] ;
    output \Add_add_temp[5] ;
    output \Add_add_temp[4] ;
    output \Error_sub_temp[30] ;
    output n31;
    input n19765;
    input n14355;
    input \qCurrent[3] ;
    input \qCurrent[4] ;
    input \qCurrent[5] ;
    input \qCurrent[6] ;
    input \qCurrent[7] ;
    input \qCurrent[8] ;
    input \qCurrent[9] ;
    input \qCurrent[10] ;
    input \qCurrent[11] ;
    input \qCurrent[12] ;
    input \qCurrent[13] ;
    input \qCurrent[14] ;
    input \qCurrent[15] ;
    input \qCurrent[16] ;
    input \qCurrent[17] ;
    input \qCurrent[18] ;
    input \qCurrent[19] ;
    input \qCurrent[20] ;
    input \qCurrent[21] ;
    input \qCurrent[22] ;
    input \qCurrent[23] ;
    input \qCurrent[24] ;
    input \qCurrent[25] ;
    input \qCurrent[26] ;
    input \qCurrent[27] ;
    input \qCurrent[28] ;
    input \qCurrent[29] ;
    input \qCurrent[30] ;
    input \qCurrent[31] ;
    input n142;
    output Saturate_out1_31__N_267;
    output Saturate_out1_31__N_266;
    input [15:0]Look_Up_Table_out1_1;
    output n579;
    output n17;
    output n267;
    output n120;
    output n14;
    output n414;
    output n11;
    output n19604;
    output n789;
    output n785;
    output n781;
    output n8;
    output n777;
    output n19351;
    output n773;
    output n769;
    output n765;
    output n270;
    output n123;
    output n761;
    output n757;
    output n417;
    output n753;
    output n749;
    output n745;
    output n741;
    output n737;
    output n489;
    output n489_adj_25;
    output n342;
    output n342_adj_26;
    output n246;
    output n288;
    output n285;
    output n282;
    output n279;
    output n276;
    output n273;
    output n258;
    output n255;
    output n252;
    output n261;
    output n249;
    output n44;
    output n126;
    output n420;
    output n129;
    output n423;
    output n41;
    output n86;
    output n89;
    output n86_adj_27;
    output n83;
    output n80;
    output n19702;
    output n77;
    output n74;
    output n38;
    output n71;
    output n68;
    output n65;
    output n62;
    output n59;
    output n56;
    output n50;
    output n53;
    output n92;
    output n244;
    output n35;
    output n195;
    output n114;
    output n108;
    output n102;
    output n99;
    output \Product2_mul_temp[2] ;
    output n141_adj_28;
    output n105;
    output n138;
    output n135;
    output n132;
    output n111;
    output n32;
    output n538;
    output n29;
    output n426;
    output n685;
    output n402;
    output n429;
    output n432;
    output n26;
    output n391;
    output n23;
    output n391_adj_29;
    output n576;
    output n576_adj_30;
    output n573;
    output n570;
    output n567;
    output n564;
    output n405;
    output n628;
    output n625;
    output n622;
    output n435;
    output n619;
    output n616;
    output n613;
    output n610;
    output n607;
    output n601;
    output n561;
    output n598;
    output n595;
    output n592;
    output n589;
    output n604;
    output n631;
    output n558;
    output n20;
    output n264;
    output n117;
    output n411;
    output n587;
    output n587_adj_31;
    output n582;
    output n393;
    output n408;
    output n555;
    output n552;
    output n549;
    output n396;
    output n399;
    output n546;
    output n543;
    output n540;
    
    wire [14:0]n841;
    wire [14:0]n842;
    
    wire n773_c, n17667, n775, n126_c, n17666;
    wire [31:0]currentControlITerm;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(59[21:40])
    
    wire n796, n17665;
    wire [31:0]preSatVoltage;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(55[22:35])
    
    wire n20174, n20858, n20870, n19884, n27, n20590, n18, n20586, 
        n20588, n20596, n20594, n20612, n20602, n20614, n20604, 
        n21, n20618, n20608, n20620, Not_Equal_relop1_N_201;
    wire [32:0]Error_sub_temp;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(44[22:36])
    wire [31:0]Proportional_Gain_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(46[22:48])
    
    wire n102_c, n737_c, n105_c, n17664, n741_c, n108_c, n745_c, 
        n111_c, n749_c, n17663, n114_c, n753_c, n117_c, n757_c, 
        n120_c, n761_c, n123_c, n765_c, n769_c, n129_c, n132_c, 
        n777_c, n135_c, n781_c, n138_c, n785_c, n789_c, n17662, 
        n17661;
    wire [14:0]n846;
    
    wire n18382, n795, n18381, n18380, n18379, n18378, n18377, 
        n18376, n18375, n18374, n18373, n18372, n18371, n18370, 
        n18369;
    wire [14:0]n845;
    
    wire n18367, n791, n18366, n18365, n18364, n18363, n18362, 
        n18361, n18360, n18359, n18358, n18357, n18356, n18355, 
        n18354;
    wire [14:0]n844;
    
    wire n18352, n787, n18351, n18350, n18349, n18348, n18347, 
        n18346, n18345, n18344, n18343, n18342, n18341, n18340, 
        n18339;
    wire [14:0]n843;
    
    wire n18337, n783, n18336, n18335, n18334, n18333, n18332, 
        n18331, n18330, n18329, n18328, n18327, n18326, n18325, 
        n18324;
    wire [14:0]n842_adj_806;
    
    wire n18322, n779, n18321, n18320, n18319, n18318, n18317, 
        n18316, n18315, n18314, n18313, n18312, n18311, n18310, 
        n18309;
    wire [14:0]n841_adj_807;
    
    wire n18307, n775_adj_590, n18306, n18305, n18304, n18303, n18302, 
        n18301, n18300, n18299, n18298, n18297, n18296, n18295, 
        n18294;
    wire [14:0]n840;
    
    wire n18292, n771, n18291, n18290, n18289, n18288, n18287, 
        n18286, n18285, n18284, n18283, n18282, n18281, n18280, 
        n18279;
    wire [14:0]n839;
    
    wire n18277, n767, n18276, n18275, n18274, n18273, n18272, 
        n18271, n18270, n18269, n18268, n18267, n18266, n18265, 
        n18264;
    wire [14:0]n838;
    
    wire n18262, n763, n18261, n18260, n18259, n18258, n18257, 
        n18256, n18255, n18254, n18253, n18252, n18251, n18250, 
        n18249;
    wire [14:0]n837;
    
    wire n18247, n759, n18246, n18245, n18244, n18243, n18242, 
        n18241, n18240, n18239, n18238, n18237, n18236, n18235, 
        n18234;
    wire [14:0]n836;
    
    wire n18232, n755, n18231, n18230, n18229, n18228, n18227, 
        n18226, n18225, n18224, n18223, n18222, n18221, n18220, 
        n18219;
    wire [14:0]n835;
    
    wire n18217, n751, n18216, n18215, n18214, n18213, n18212, 
        n18211, n18210, n18209, n18208, n18207, n18206, n18205, 
        n18204;
    wire [14:0]n834;
    
    wire n18202, n747, n18201, n18200, n18199, n18198, n18197, 
        n18196, n18195, n18194, n18193, n18192, n18191, n18190, 
        n18189;
    wire [14:0]n833;
    
    wire n18187, n743, n18186;
    wire [31:0]Switch_out1;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(58[22:33])
    
    wire n18185, n18184, n18183, n18182, n18181, n18180, n18179, 
        n18178, n18177, n18176, n18175, n18174, n18159, n18158, 
        n18157, n18156, n18155, n18154, n18153, n18152, n18151, 
        n18150, n18149, n18148, n18147, n18146, n8356, n18145, 
        n18144;
    wire [14:0]n832;
    wire [14:0]n840_adj_808;
    
    wire n18120, n771_adj_598, n18119, n18118, n18117, n18116, n18115, 
        n18114, n18113, n18112, n18111, n18110, n18109, n18108, 
        n18107;
    wire [14:0]n839_adj_809;
    
    wire n18105, n767_adj_620, n18104, n18103, n18102, n18101, n18100, 
        n18099, n18098, n18097, n18096, n18095, n18094, n18093, 
        n18092;
    wire [14:0]n838_adj_810;
    
    wire n18090, n763_adj_636, n18089, n18088, n18087, n18086, n18085, 
        n18084, n18083, n18082, n18081, n18080, n18079, n18078, 
        n18077;
    wire [14:0]n837_adj_811;
    
    wire n18075, n759_adj_652, n18074, n18073, n18072, n18071, n18070, 
        n18069, n18068, n18067, n18066, n18065, n18064, n18063, 
        n18062;
    wire [14:0]n836_adj_812;
    
    wire n18060, n755_adj_668, n18059, n18058, n18057, n18056, n18055, 
        n18054, n18053, n18052, n18051, n18050, n18049, n18048, 
        n18047;
    wire [14:0]n835_adj_813;
    
    wire n18045, n751_adj_684, n18044, n18043, n18042, n18041, n18040, 
        n18039, n18038, n18037, n18036, n18035, n18034, n18033, 
        n18032;
    wire [14:0]n834_adj_814;
    
    wire n18030, n747_adj_700, n18029, n18028, n18027, n18026, n18025, 
        n18024, n18023, n18022, n18021, n18020, n18019, n18018, 
        n18017;
    wire [14:0]n833_adj_815;
    
    wire n18015, n743_adj_716, n18014, n18013, n18012, n18011, n18010, 
        n18009, n18008, n18007, n18006, n18005, n18004, n18003, 
        n18002;
    wire [14:0]n832_adj_816;
    
    wire n18000, n739, n17999, n17998, n17997, n17996, n17995, 
        n17994, n17993, n17992, n17991, n17990, n17989, n17988, 
        n17987;
    wire [14:0]n844_adj_817;
    wire [14:0]n845_adj_818;
    
    wire n17978, n787_adj_721, n17977, n17976, n17975, n17974, n17973, 
        n17972, n791_adj_732, n17971, n17970, n783_adj_734, n17969;
    wire [14:0]n843_adj_819;
    
    wire n779_adj_736, n17968, n17967, n17966, n17965, n17964, n17963, 
        n17962, n17961, n17960, n17959, n17958, n17957, n17734, 
        n17733, n17732, n17731, n17660, n17659, n17730, n17865, 
        n17864, n17863, n17862;
    wire [31:0]Saturate_out1;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(64[22:35])
    
    wire n15943, n15942, n15941, n17861, n15940, n15939, n17860, 
        n17859, n15938, n15937, n15936, n15935, n15934, n15933, 
        n15932, n15931, n15930, n15929, n15928, n15927, n15926, 
        n15925, n15924, n15923, n15922, n15921, n15920, n15919, 
        n15918, n15917, n15916, n15915, n15914, n15913;
    wire [31:0]Voltage_1;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(56[22:31])
    
    wire n15912, n15911, n15910, n15909, n15908, n15907, n15906, 
        n15905, n15904, n15903, n15902, n15901, n15900, n15899, 
        n15898, n15897, n15896, n15895, n15894, n15893, n15892, 
        n15891, n15890, n15889, n15888, n15887, n15886, n15885, 
        n15884, n15883, n17858, n17857, n17658, n17856, n17729, 
        n17657, n17728, n17656, n17727;
    wire [29:0]n1;
    
    wire n15747, n15746, n15745, n15744, n15743, n15742, n15741, 
        n15740, n15739, n15738, n15737, n15736, n15735, n15734, 
        n15733, n15732, n15731, n15730, n15729, n15728, n15727, 
        n15726, n15725, n15724, n15723, n15722, n15721, n15720, 
        n10_adj_755, n14_adj_756, n4_adj_757, n18_adj_758, n19841, 
        n26_adj_759, n7_adj_760, n4_adj_761, n20722, n19761, n20704, 
        n15200, n20680, n19733, n20660, n20654, n20640, n19308, 
        n19755, n20718, n22_adj_762, n20694, n19729, n20676, n20664, 
        n20650, n58, n6_adj_763;
    
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_14_lut (.I0(GND_net), .I1(n842[9]), 
            .I2(n773_c), .I3(n17667), .O(n841[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_14 (.CI(n17667), .I0(n842[9]), 
            .I1(n773_c), .CO(n775));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_13_lut (.I0(GND_net), .I1(n842[9]), 
            .I2(n126_c), .I3(n17666), .O(n841[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_13 (.CI(n17666), .I0(n842[9]), 
            .I1(n126_c), .CO(n17667));
    SB_DFF currentControlITerm_i30 (.Q(currentControlITerm[30]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14381));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 paramCurrentControlP_15__I_0_i542_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(\Error_sub_temp[31] ), .I2(GND_net), .I3(GND_net), .O(n796));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i542_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_12_lut (.I0(GND_net), .I1(n842[9]), 
            .I2(n126_c), .I3(n17665), .O(n841[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_12 (.CI(n17665), .I0(n842[9]), 
            .I1(n126_c), .CO(n17666));
    SB_LUT4 i15877_4_lut (.I0(preSatVoltage[4]), .I1(preSatVoltage[3]), 
            .I2(preSatVoltage[2]), .I3(n20174), .O(n20858));
    defparam i15877_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15889_4_lut (.I0(preSatVoltage[7]), .I1(preSatVoltage[6]), 
            .I2(preSatVoltage[5]), .I3(n20858), .O(n20870));
    defparam i15889_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(\preSatVoltage[10] ), .I1(preSatVoltage[9]), .I2(preSatVoltage[8]), 
            .I3(n20870), .O(n19884));
    defparam i1_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 equal_13244_i27_3_lut (.I0(preSatVoltage[26]), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(n27));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam equal_13244_i27_3_lut.LUT_INIT = 16'ha4a4;
    SB_LUT4 i1_4_lut_adj_260 (.I0(preSatVoltage[28]), .I1(preSatVoltage[29]), 
            .I2(Out_31__N_333), .I3(Out_31__N_332), .O(n20590));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_260.LUT_INIT = 16'hee70;
    SB_LUT4 equal_13244_i18_2_lut (.I0(preSatVoltage[17]), .I1(\qVoltage[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam equal_13244_i18_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_261 (.I0(preSatVoltage[27]), .I1(n19884), .I2(Out_31__N_333), 
            .I3(Out_31__N_332), .O(n20586));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_261.LUT_INIT = 16'hbb70;
    SB_LUT4 i1_4_lut_adj_262 (.I0(preSatVoltage[30]), .I1(preSatVoltage[25]), 
            .I2(Out_31__N_333), .I3(Out_31__N_332), .O(n20588));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_262.LUT_INIT = 16'hee70;
    SB_LUT4 i1_3_lut (.I0(n20588), .I1(preSatVoltage[14]), .I2(\qVoltage[5] ), 
            .I3(GND_net), .O(n20596));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i1_4_lut_adj_263 (.I0(preSatVoltage[11]), .I1(preSatVoltage[21]), 
            .I2(\qVoltage[2] ), .I3(\qVoltage[12] ), .O(n20594));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_263.LUT_INIT = 16'h7bde;
    SB_DFF currentControlITerm_i29 (.Q(currentControlITerm[29]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14380));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 i1_4_lut_adj_264 (.I0(\preSatVoltage[23] ), .I1(preSatVoltage[18]), 
            .I2(\qVoltage[14] ), .I3(\qVoltage[9] ), .O(n20612));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_264.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_265 (.I0(n20586), .I1(n18), .I2(n20590), .I3(n27), 
            .O(n20602));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_265.LUT_INIT = 16'hfffe;
    SB_DFF currentControlITerm_i28 (.Q(currentControlITerm[28]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14379));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 i1_4_lut_adj_266 (.I0(\preSatVoltage[13] ), .I1(\preSatVoltage[12] ), 
            .I2(\qVoltage[4] ), .I3(\qVoltage[3] ), .O(n20614));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_266.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_267 (.I0(n20594), .I1(n20596), .I2(preSatVoltage[24]), 
            .I3(\qVoltage[15] ), .O(n20604));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_267.LUT_INIT = 16'heffe;
    SB_DFF currentControlITerm_i27 (.Q(currentControlITerm[27]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14378));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i26 (.Q(currentControlITerm[26]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14377));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i25 (.Q(currentControlITerm[25]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14376));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i24 (.Q(currentControlITerm[24]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14375));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i23 (.Q(currentControlITerm[23]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14374));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 i1_4_lut_adj_268 (.I0(preSatVoltage[15]), .I1(n20612), .I2(n21), 
            .I3(\qVoltage[6] ), .O(n20618));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_268.LUT_INIT = 16'hfdfe;
    SB_DFF currentControlITerm_i22 (.Q(currentControlITerm[22]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14373));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 i1_4_lut_adj_269 (.I0(\preSatVoltage[22] ), .I1(\preSatVoltage[19] ), 
            .I2(\qVoltage[13] ), .I3(\qVoltage[10] ), .O(n20608));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_269.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_270 (.I0(n20614), .I1(preSatVoltage[16]), .I2(n20602), 
            .I3(\qVoltage[7] ), .O(n20620));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_270.LUT_INIT = 16'hfbfe;
    SB_LUT4 equal_13244_i62_4_lut (.I0(n20620), .I1(n20608), .I2(n20618), 
            .I3(n20604), .O(Not_Equal_relop1_N_201));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam equal_13244_i62_4_lut.LUT_INIT = 16'h0001;
    SB_DFF currentControlITerm_i3 (.Q(currentControlITerm[3]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14354));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i21 (.Q(currentControlITerm[21]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14372));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i20 (.Q(currentControlITerm[20]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14371));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i19 (.Q(currentControlITerm[19]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14370));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i18 (.Q(currentControlITerm[18]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14369));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i2 (.Q(currentControlITerm[2]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14353));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i17 (.Q(currentControlITerm[17]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14368));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i16 (.Q(currentControlITerm[16]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14367));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i15 (.Q(currentControlITerm[15]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14366));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i14 (.Q(currentControlITerm[14]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14365));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i13 (.Q(currentControlITerm[13]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14364));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i12 (.Q(currentControlITerm[12]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14363));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i11 (.Q(currentControlITerm[11]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14362));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i10 (.Q(currentControlITerm[10]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14361));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i9 (.Q(currentControlITerm[9]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14360));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i8 (.Q(currentControlITerm[8]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14359));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i1 (.Q(currentControlITerm[1]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14352));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 paramCurrentControlP_15__I_0_i35_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[16]), .I2(GND_net), .I3(GND_net), .O(Proportional_Gain_mul_temp[0]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i35_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i37_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[17]), .I2(GND_net), .I3(GND_net), .O(n102_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i37_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i498_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[16]), .I2(GND_net), .I3(GND_net), .O(n737_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i498_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i39_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[18]), .I2(GND_net), .I3(GND_net), .O(n105_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i39_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_11_lut (.I0(GND_net), .I1(n842[8]), 
            .I2(n126_c), .I3(n17664), .O(n841[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_i501_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[17]), .I2(GND_net), .I3(GND_net), .O(n741_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i501_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_11 (.CI(n17664), .I0(n842[8]), 
            .I1(n126_c), .CO(n17665));
    SB_LUT4 paramCurrentControlP_15__I_0_i41_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[19]), .I2(GND_net), .I3(GND_net), .O(n108_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i41_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i504_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[18]), .I2(GND_net), .I3(GND_net), .O(n745_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i504_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i43_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[20]), .I2(GND_net), .I3(GND_net), .O(n111_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i43_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i507_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[19]), .I2(GND_net), .I3(GND_net), .O(n749_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i507_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_10_lut (.I0(GND_net), .I1(n842[7]), 
            .I2(n126_c), .I3(n17663), .O(n841[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_i45_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[21]), .I2(GND_net), .I3(GND_net), .O(n114_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i45_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i510_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[20]), .I2(GND_net), .I3(GND_net), .O(n753_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i510_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i47_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[22]), .I2(GND_net), .I3(GND_net), .O(n117_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i47_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i513_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[21]), .I2(GND_net), .I3(GND_net), .O(n757_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i513_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i49_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[23]), .I2(GND_net), .I3(GND_net), .O(n120_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i49_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_10 (.CI(n17663), .I0(n842[7]), 
            .I1(n126_c), .CO(n17664));
    SB_LUT4 paramCurrentControlP_15__I_0_i516_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[22]), .I2(GND_net), .I3(GND_net), .O(n761_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i516_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i51_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[24]), .I2(GND_net), .I3(GND_net), .O(n123_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i51_2_lut.LUT_INIT = 16'h8888;
    SB_DFF currentControlITerm_i7 (.Q(preSatVoltage[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14358));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 paramCurrentControlP_15__I_0_i519_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[23]), .I2(GND_net), .I3(GND_net), .O(n765_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i519_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i522_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[24]), .I2(GND_net), .I3(GND_net), .O(n769_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i522_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i55_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[26]), .I2(GND_net), .I3(GND_net), .O(n129_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i57_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[27]), .I2(GND_net), .I3(GND_net), .O(n132_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i528_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[26]), .I2(GND_net), .I3(GND_net), .O(n777_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i528_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i59_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[28]), .I2(GND_net), .I3(GND_net), .O(n135_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i531_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[27]), .I2(GND_net), .I3(GND_net), .O(n781_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i531_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i61_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[29]), .I2(GND_net), .I3(GND_net), .O(n138_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i534_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[28]), .I2(GND_net), .I3(GND_net), .O(n785_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i534_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i537_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[29]), .I2(GND_net), .I3(GND_net), .O(n789_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i537_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_9_lut (.I0(GND_net), .I1(n842[6]), 
            .I2(n126_c), .I3(n17662), .O(n841[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_i66_2_lut (.I0(\Amp25_out1[14] ), 
            .I1(\Error_sub_temp[31] ), .I2(GND_net), .I3(GND_net), .O(n146));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i66_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_9 (.CI(n17662), .I0(n842[6]), 
            .I1(n126_c), .CO(n17663));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_8_lut (.I0(GND_net), .I1(n842[5]), 
            .I2(n126_c), .I3(n17661), .O(n841[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF currentControlITerm_i6 (.Q(currentControlITerm[6]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14357));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i5 (.Q(currentControlITerm[5]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14356));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 Error_sub_temp_31__I_0_add_575_16_lut (.I0(GND_net), .I1(n793), 
            .I2(n146), .I3(n18382), .O(n846[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_16 (.CI(n18382), .I0(n793), 
            .I1(n146), .CO(n795));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_15_lut (.I0(GND_net), .I1(n789_c), 
            .I2(n141), .I3(n18381), .O(n846[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_15 (.CI(n18381), .I0(n789_c), 
            .I1(n141), .CO(n18382));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_14_lut (.I0(GND_net), .I1(n785_c), 
            .I2(n138_c), .I3(n18380), .O(n846[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_14 (.CI(n18380), .I0(n785_c), 
            .I1(n138_c), .CO(n18381));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_13_lut (.I0(GND_net), .I1(n781_c), 
            .I2(n135_c), .I3(n18379), .O(n846[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_13 (.CI(n18379), .I0(n781_c), 
            .I1(n135_c), .CO(n18380));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_12_lut (.I0(GND_net), .I1(n777_c), 
            .I2(n132_c), .I3(n18378), .O(n846[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_12 (.CI(n18378), .I0(n777_c), 
            .I1(n132_c), .CO(n18379));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_11_lut (.I0(GND_net), .I1(n773_c), 
            .I2(n129_c), .I3(n18377), .O(n846[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_11 (.CI(n18377), .I0(n773_c), 
            .I1(n129_c), .CO(n18378));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_10_lut (.I0(GND_net), .I1(n769_c), 
            .I2(n126_c), .I3(n18376), .O(n846[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_10 (.CI(n18376), .I0(n769_c), 
            .I1(n126_c), .CO(n18377));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_9_lut (.I0(GND_net), .I1(n765_c), 
            .I2(n123_c), .I3(n18375), .O(n846[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_9 (.CI(n18375), .I0(n765_c), 
            .I1(n123_c), .CO(n18376));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_8_lut (.I0(GND_net), .I1(n761_c), 
            .I2(n120_c), .I3(n18374), .O(n846[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_8 (.CI(n18374), .I0(n761_c), 
            .I1(n120_c), .CO(n18375));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_7_lut (.I0(GND_net), .I1(n757_c), 
            .I2(n117_c), .I3(n18373), .O(n846[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_7 (.CI(n18373), .I0(n757_c), 
            .I1(n117_c), .CO(n18374));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_6_lut (.I0(GND_net), .I1(n753_c), 
            .I2(n114_c), .I3(n18372), .O(n846[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_6 (.CI(n18372), .I0(n753_c), 
            .I1(n114_c), .CO(n18373));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_5_lut (.I0(GND_net), .I1(n749_c), 
            .I2(n111_c), .I3(n18371), .O(n846[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_5 (.CI(n18371), .I0(n749_c), 
            .I1(n111_c), .CO(n18372));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_4_lut (.I0(GND_net), .I1(n745_c), 
            .I2(n108_c), .I3(n18370), .O(n846[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_4 (.CI(n18370), .I0(n745_c), 
            .I1(n108_c), .CO(n18371));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_3_lut (.I0(GND_net), .I1(n741_c), 
            .I2(n105_c), .I3(n18369), .O(n846[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_3 (.CI(n18369), .I0(n741_c), 
            .I1(n105_c), .CO(n18370));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_2_lut (.I0(GND_net), .I1(n737_c), 
            .I2(n102_c), .I3(GND_net), .O(n846[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_2 (.CI(GND_net), .I0(n737_c), 
            .I1(n102_c), .CO(n18369));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_16_lut (.I0(GND_net), .I1(n846[13]), 
            .I2(n146), .I3(n18367), .O(n845[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_16 (.CI(n18367), .I0(n846[13]), 
            .I1(n146), .CO(n791));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_15_lut (.I0(GND_net), .I1(n846[12]), 
            .I2(n141), .I3(n18366), .O(n845[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_15 (.CI(n18366), .I0(n846[12]), 
            .I1(n141), .CO(n18367));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_14_lut (.I0(GND_net), .I1(n846[11]), 
            .I2(n138_c), .I3(n18365), .O(n845[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_14 (.CI(n18365), .I0(n846[11]), 
            .I1(n138_c), .CO(n18366));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_13_lut (.I0(GND_net), .I1(n846[10]), 
            .I2(n135_c), .I3(n18364), .O(n845[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_13 (.CI(n18364), .I0(n846[10]), 
            .I1(n135_c), .CO(n18365));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_12_lut (.I0(GND_net), .I1(n846[9]), 
            .I2(n132_c), .I3(n18363), .O(n845[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_12 (.CI(n18363), .I0(n846[9]), 
            .I1(n132_c), .CO(n18364));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_11_lut (.I0(GND_net), .I1(n846[8]), 
            .I2(n129_c), .I3(n18362), .O(n845[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_11 (.CI(n18362), .I0(n846[8]), 
            .I1(n129_c), .CO(n18363));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_10_lut (.I0(GND_net), .I1(n846[7]), 
            .I2(n126_c), .I3(n18361), .O(n845[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_10 (.CI(n18361), .I0(n846[7]), 
            .I1(n126_c), .CO(n18362));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_9_lut (.I0(GND_net), .I1(n846[6]), 
            .I2(n123_c), .I3(n18360), .O(n845[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_9 (.CI(n18360), .I0(n846[6]), 
            .I1(n123_c), .CO(n18361));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_8_lut (.I0(GND_net), .I1(n846[5]), 
            .I2(n120_c), .I3(n18359), .O(n845[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_8 (.CI(n18359), .I0(n846[5]), 
            .I1(n120_c), .CO(n18360));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_7_lut (.I0(GND_net), .I1(n846[4]), 
            .I2(n117_c), .I3(n18358), .O(n845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_7 (.CI(n18358), .I0(n846[4]), 
            .I1(n117_c), .CO(n18359));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_6_lut (.I0(GND_net), .I1(n846[3]), 
            .I2(n114_c), .I3(n18357), .O(n845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_6 (.CI(n18357), .I0(n846[3]), 
            .I1(n114_c), .CO(n18358));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_5_lut (.I0(GND_net), .I1(n846[2]), 
            .I2(n111_c), .I3(n18356), .O(n845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_5 (.CI(n18356), .I0(n846[2]), 
            .I1(n111_c), .CO(n18357));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_4_lut (.I0(GND_net), .I1(n846[1]), 
            .I2(n108_c), .I3(n18355), .O(n845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_4 (.CI(n18355), .I0(n846[1]), 
            .I1(n108_c), .CO(n18356));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_3_lut (.I0(GND_net), .I1(n846[0]), 
            .I2(n105_c), .I3(n18354), .O(n845[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_3 (.CI(n18354), .I0(n846[0]), 
            .I1(n105_c), .CO(n18355));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n845[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18354));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_16_lut (.I0(GND_net), .I1(n845[13]), 
            .I2(n146), .I3(n18352), .O(n844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_16 (.CI(n18352), .I0(n845[13]), 
            .I1(n146), .CO(n787));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_15_lut (.I0(GND_net), .I1(n845[12]), 
            .I2(n141), .I3(n18351), .O(n844[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_15 (.CI(n18351), .I0(n845[12]), 
            .I1(n141), .CO(n18352));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_14_lut (.I0(GND_net), .I1(n845[11]), 
            .I2(n138_c), .I3(n18350), .O(n844[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_14 (.CI(n18350), .I0(n845[11]), 
            .I1(n138_c), .CO(n18351));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_13_lut (.I0(GND_net), .I1(n845[10]), 
            .I2(n135_c), .I3(n18349), .O(n844[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_13 (.CI(n18349), .I0(n845[10]), 
            .I1(n135_c), .CO(n18350));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_12_lut (.I0(GND_net), .I1(n845[9]), 
            .I2(n132_c), .I3(n18348), .O(n844[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_12 (.CI(n18348), .I0(n845[9]), 
            .I1(n132_c), .CO(n18349));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_11_lut (.I0(GND_net), .I1(n845[8]), 
            .I2(n129_c), .I3(n18347), .O(n844[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_11 (.CI(n18347), .I0(n845[8]), 
            .I1(n129_c), .CO(n18348));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_10_lut (.I0(GND_net), .I1(n845[7]), 
            .I2(n126_c), .I3(n18346), .O(n844[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_10 (.CI(n18346), .I0(n845[7]), 
            .I1(n126_c), .CO(n18347));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_9_lut (.I0(GND_net), .I1(n845[6]), 
            .I2(n123_c), .I3(n18345), .O(n844[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_9 (.CI(n18345), .I0(n845[6]), 
            .I1(n123_c), .CO(n18346));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_8_lut (.I0(GND_net), .I1(n845[5]), 
            .I2(n120_c), .I3(n18344), .O(n844[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_8 (.CI(n18344), .I0(n845[5]), 
            .I1(n120_c), .CO(n18345));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_7_lut (.I0(GND_net), .I1(n845[4]), 
            .I2(n117_c), .I3(n18343), .O(n844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_7 (.CI(n18343), .I0(n845[4]), 
            .I1(n117_c), .CO(n18344));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_6_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n114_c), .I3(n18342), .O(n844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_6 (.CI(n18342), .I0(n845[3]), 
            .I1(n114_c), .CO(n18343));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_5_lut (.I0(GND_net), .I1(n845[2]), 
            .I2(n111_c), .I3(n18341), .O(n844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_5 (.CI(n18341), .I0(n845[2]), 
            .I1(n111_c), .CO(n18342));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_4_lut (.I0(GND_net), .I1(n845[1]), 
            .I2(n108_c), .I3(n18340), .O(n844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_4 (.CI(n18340), .I0(n845[1]), 
            .I1(n108_c), .CO(n18341));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_3_lut (.I0(GND_net), .I1(n845[0]), 
            .I2(n105_c), .I3(n18339), .O(n844[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_3 (.CI(n18339), .I0(n845[0]), 
            .I1(n105_c), .CO(n18340));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n844[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18339));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_16_lut (.I0(GND_net), .I1(n844[13]), 
            .I2(n146), .I3(n18337), .O(n843[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_16 (.CI(n18337), .I0(n844[13]), 
            .I1(n146), .CO(n783));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_15_lut (.I0(GND_net), .I1(n844[12]), 
            .I2(n141), .I3(n18336), .O(n843[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_15 (.CI(n18336), .I0(n844[12]), 
            .I1(n141), .CO(n18337));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_14_lut (.I0(GND_net), .I1(n844[11]), 
            .I2(n138_c), .I3(n18335), .O(n843[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_14 (.CI(n18335), .I0(n844[11]), 
            .I1(n138_c), .CO(n18336));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_13_lut (.I0(GND_net), .I1(n844[10]), 
            .I2(n135_c), .I3(n18334), .O(n843[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_13 (.CI(n18334), .I0(n844[10]), 
            .I1(n135_c), .CO(n18335));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_12_lut (.I0(GND_net), .I1(n844[9]), 
            .I2(n132_c), .I3(n18333), .O(n843[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_12 (.CI(n18333), .I0(n844[9]), 
            .I1(n132_c), .CO(n18334));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_11_lut (.I0(GND_net), .I1(n844[8]), 
            .I2(n129_c), .I3(n18332), .O(n843[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_11 (.CI(n18332), .I0(n844[8]), 
            .I1(n129_c), .CO(n18333));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_10_lut (.I0(GND_net), .I1(n844[7]), 
            .I2(n126_c), .I3(n18331), .O(n843[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_10 (.CI(n18331), .I0(n844[7]), 
            .I1(n126_c), .CO(n18332));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_9_lut (.I0(GND_net), .I1(n844[6]), 
            .I2(n123_c), .I3(n18330), .O(n843[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_9 (.CI(n18330), .I0(n844[6]), 
            .I1(n123_c), .CO(n18331));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_8_lut (.I0(GND_net), .I1(n844[5]), 
            .I2(n120_c), .I3(n18329), .O(n843[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_8 (.CI(n18329), .I0(n844[5]), 
            .I1(n120_c), .CO(n18330));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_7_lut (.I0(GND_net), .I1(n844[4]), 
            .I2(n117_c), .I3(n18328), .O(n843[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_7 (.CI(n18328), .I0(n844[4]), 
            .I1(n117_c), .CO(n18329));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_6_lut (.I0(GND_net), .I1(n844[3]), 
            .I2(n114_c), .I3(n18327), .O(n843[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_6 (.CI(n18327), .I0(n844[3]), 
            .I1(n114_c), .CO(n18328));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_5_lut (.I0(GND_net), .I1(n844[2]), 
            .I2(n111_c), .I3(n18326), .O(n843[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_5 (.CI(n18326), .I0(n844[2]), 
            .I1(n111_c), .CO(n18327));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_4_lut (.I0(GND_net), .I1(n844[1]), 
            .I2(n108_c), .I3(n18325), .O(n843[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_4 (.CI(n18325), .I0(n844[1]), 
            .I1(n108_c), .CO(n18326));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_3_lut (.I0(GND_net), .I1(n844[0]), 
            .I2(n105_c), .I3(n18324), .O(n843[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_3 (.CI(n18324), .I0(n844[0]), 
            .I1(n105_c), .CO(n18325));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n843[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18324));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_16_lut (.I0(GND_net), .I1(n843[13]), 
            .I2(n146), .I3(n18322), .O(n842_adj_806[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_16 (.CI(n18322), .I0(n843[13]), 
            .I1(n146), .CO(n779));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_15_lut (.I0(GND_net), .I1(n843[12]), 
            .I2(n141), .I3(n18321), .O(n842_adj_806[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_15 (.CI(n18321), .I0(n843[12]), 
            .I1(n141), .CO(n18322));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_14_lut (.I0(GND_net), .I1(n843[11]), 
            .I2(n138_c), .I3(n18320), .O(n842_adj_806[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_14 (.CI(n18320), .I0(n843[11]), 
            .I1(n138_c), .CO(n18321));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_13_lut (.I0(GND_net), .I1(n843[10]), 
            .I2(n135_c), .I3(n18319), .O(n842_adj_806[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_13 (.CI(n18319), .I0(n843[10]), 
            .I1(n135_c), .CO(n18320));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_12_lut (.I0(GND_net), .I1(n843[9]), 
            .I2(n132_c), .I3(n18318), .O(n842_adj_806[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_12 (.CI(n18318), .I0(n843[9]), 
            .I1(n132_c), .CO(n18319));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_11_lut (.I0(GND_net), .I1(n843[8]), 
            .I2(n129_c), .I3(n18317), .O(n842_adj_806[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_11 (.CI(n18317), .I0(n843[8]), 
            .I1(n129_c), .CO(n18318));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_10_lut (.I0(GND_net), .I1(n843[7]), 
            .I2(n126_c), .I3(n18316), .O(n842_adj_806[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_10 (.CI(n18316), .I0(n843[7]), 
            .I1(n126_c), .CO(n18317));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_9_lut (.I0(GND_net), .I1(n843[6]), 
            .I2(n123_c), .I3(n18315), .O(n842_adj_806[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_9 (.CI(n18315), .I0(n843[6]), 
            .I1(n123_c), .CO(n18316));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_8_lut (.I0(GND_net), .I1(n843[5]), 
            .I2(n120_c), .I3(n18314), .O(n842_adj_806[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_8 (.CI(n18314), .I0(n843[5]), 
            .I1(n120_c), .CO(n18315));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_7_lut (.I0(GND_net), .I1(n843[4]), 
            .I2(n117_c), .I3(n18313), .O(n842_adj_806[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_7 (.CI(n18313), .I0(n843[4]), 
            .I1(n117_c), .CO(n18314));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_6_lut (.I0(GND_net), .I1(n843[3]), 
            .I2(n114_c), .I3(n18312), .O(n842_adj_806[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_6 (.CI(n18312), .I0(n843[3]), 
            .I1(n114_c), .CO(n18313));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_5_lut (.I0(GND_net), .I1(n843[2]), 
            .I2(n111_c), .I3(n18311), .O(n842_adj_806[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_5 (.CI(n18311), .I0(n843[2]), 
            .I1(n111_c), .CO(n18312));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_4_lut (.I0(GND_net), .I1(n843[1]), 
            .I2(n108_c), .I3(n18310), .O(n842_adj_806[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_4 (.CI(n18310), .I0(n843[1]), 
            .I1(n108_c), .CO(n18311));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_3_lut (.I0(GND_net), .I1(n843[0]), 
            .I2(n105_c), .I3(n18309), .O(n842_adj_806[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_3 (.CI(n18309), .I0(n843[0]), 
            .I1(n105_c), .CO(n18310));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n842_adj_806[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18309));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_16_lut (.I0(GND_net), .I1(n842_adj_806[13]), 
            .I2(n146), .I3(n18307), .O(n841_adj_807[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_16 (.CI(n18307), .I0(n842_adj_806[13]), 
            .I1(n146), .CO(n775_adj_590));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_15_lut (.I0(GND_net), .I1(n842_adj_806[12]), 
            .I2(n141), .I3(n18306), .O(n841_adj_807[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_15 (.CI(n18306), .I0(n842_adj_806[12]), 
            .I1(n141), .CO(n18307));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_14_lut (.I0(GND_net), .I1(n842_adj_806[11]), 
            .I2(n138_c), .I3(n18305), .O(n841_adj_807[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_14 (.CI(n18305), .I0(n842_adj_806[11]), 
            .I1(n138_c), .CO(n18306));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_13_lut (.I0(GND_net), .I1(n842_adj_806[10]), 
            .I2(n135_c), .I3(n18304), .O(n841_adj_807[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_13 (.CI(n18304), .I0(n842_adj_806[10]), 
            .I1(n135_c), .CO(n18305));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_12_lut (.I0(GND_net), .I1(n842_adj_806[9]), 
            .I2(n132_c), .I3(n18303), .O(n841_adj_807[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_12 (.CI(n18303), .I0(n842_adj_806[9]), 
            .I1(n132_c), .CO(n18304));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_11_lut (.I0(GND_net), .I1(n842_adj_806[8]), 
            .I2(n129_c), .I3(n18302), .O(n841_adj_807[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_11 (.CI(n18302), .I0(n842_adj_806[8]), 
            .I1(n129_c), .CO(n18303));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_10_lut (.I0(GND_net), .I1(n842_adj_806[7]), 
            .I2(n126_c), .I3(n18301), .O(n841_adj_807[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_10 (.CI(n18301), .I0(n842_adj_806[7]), 
            .I1(n126_c), .CO(n18302));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_9_lut (.I0(GND_net), .I1(n842_adj_806[6]), 
            .I2(n123_c), .I3(n18300), .O(n841_adj_807[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_9 (.CI(n18300), .I0(n842_adj_806[6]), 
            .I1(n123_c), .CO(n18301));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_8_lut (.I0(GND_net), .I1(n842_adj_806[5]), 
            .I2(n120_c), .I3(n18299), .O(n841_adj_807[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_8 (.CI(n18299), .I0(n842_adj_806[5]), 
            .I1(n120_c), .CO(n18300));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_7_lut (.I0(GND_net), .I1(n842_adj_806[4]), 
            .I2(n117_c), .I3(n18298), .O(n841_adj_807[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_7 (.CI(n18298), .I0(n842_adj_806[4]), 
            .I1(n117_c), .CO(n18299));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_6_lut (.I0(GND_net), .I1(n842_adj_806[3]), 
            .I2(n114_c), .I3(n18297), .O(n841_adj_807[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_6 (.CI(n18297), .I0(n842_adj_806[3]), 
            .I1(n114_c), .CO(n18298));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_5_lut (.I0(GND_net), .I1(n842_adj_806[2]), 
            .I2(n111_c), .I3(n18296), .O(n841_adj_807[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_5 (.CI(n18296), .I0(n842_adj_806[2]), 
            .I1(n111_c), .CO(n18297));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_4_lut (.I0(GND_net), .I1(n842_adj_806[1]), 
            .I2(n108_c), .I3(n18295), .O(n841_adj_807[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_4 (.CI(n18295), .I0(n842_adj_806[1]), 
            .I1(n108_c), .CO(n18296));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_3_lut (.I0(GND_net), .I1(n842_adj_806[0]), 
            .I2(n105_c), .I3(n18294), .O(n841_adj_807[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_3 (.CI(n18294), .I0(n842_adj_806[0]), 
            .I1(n105_c), .CO(n18295));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n841_adj_807[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18294));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_16_lut (.I0(GND_net), .I1(n841_adj_807[13]), 
            .I2(n146), .I3(n18292), .O(n840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_16 (.CI(n18292), .I0(n841_adj_807[13]), 
            .I1(n146), .CO(n771));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_15_lut (.I0(GND_net), .I1(n841_adj_807[12]), 
            .I2(n141), .I3(n18291), .O(n840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_15 (.CI(n18291), .I0(n841_adj_807[12]), 
            .I1(n141), .CO(n18292));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_14_lut (.I0(GND_net), .I1(n841_adj_807[11]), 
            .I2(n138_c), .I3(n18290), .O(n840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_14 (.CI(n18290), .I0(n841_adj_807[11]), 
            .I1(n138_c), .CO(n18291));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_13_lut (.I0(GND_net), .I1(n841_adj_807[10]), 
            .I2(n135_c), .I3(n18289), .O(n840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_13 (.CI(n18289), .I0(n841_adj_807[10]), 
            .I1(n135_c), .CO(n18290));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_12_lut (.I0(GND_net), .I1(n841_adj_807[9]), 
            .I2(n132_c), .I3(n18288), .O(n840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_12 (.CI(n18288), .I0(n841_adj_807[9]), 
            .I1(n132_c), .CO(n18289));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_11_lut (.I0(GND_net), .I1(n841_adj_807[8]), 
            .I2(n129_c), .I3(n18287), .O(n840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_11 (.CI(n18287), .I0(n841_adj_807[8]), 
            .I1(n129_c), .CO(n18288));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_10_lut (.I0(GND_net), .I1(n841_adj_807[7]), 
            .I2(n126_c), .I3(n18286), .O(n840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_10 (.CI(n18286), .I0(n841_adj_807[7]), 
            .I1(n126_c), .CO(n18287));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_9_lut (.I0(GND_net), .I1(n841_adj_807[6]), 
            .I2(n123_c), .I3(n18285), .O(n840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_9 (.CI(n18285), .I0(n841_adj_807[6]), 
            .I1(n123_c), .CO(n18286));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_8_lut (.I0(GND_net), .I1(n841_adj_807[5]), 
            .I2(n120_c), .I3(n18284), .O(n840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_8 (.CI(n18284), .I0(n841_adj_807[5]), 
            .I1(n120_c), .CO(n18285));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_7_lut (.I0(GND_net), .I1(n841_adj_807[4]), 
            .I2(n117_c), .I3(n18283), .O(n840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_7 (.CI(n18283), .I0(n841_adj_807[4]), 
            .I1(n117_c), .CO(n18284));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_6_lut (.I0(GND_net), .I1(n841_adj_807[3]), 
            .I2(n114_c), .I3(n18282), .O(n840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_6 (.CI(n18282), .I0(n841_adj_807[3]), 
            .I1(n114_c), .CO(n18283));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_5_lut (.I0(GND_net), .I1(n841_adj_807[2]), 
            .I2(n111_c), .I3(n18281), .O(n840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_5 (.CI(n18281), .I0(n841_adj_807[2]), 
            .I1(n111_c), .CO(n18282));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_4_lut (.I0(GND_net), .I1(n841_adj_807[1]), 
            .I2(n108_c), .I3(n18280), .O(n840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_4 (.CI(n18280), .I0(n841_adj_807[1]), 
            .I1(n108_c), .CO(n18281));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_3_lut (.I0(GND_net), .I1(n841_adj_807[0]), 
            .I2(n105_c), .I3(n18279), .O(n840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_3 (.CI(n18279), .I0(n841_adj_807[0]), 
            .I1(n105_c), .CO(n18280));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18279));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_16_lut (.I0(GND_net), .I1(n840[13]), 
            .I2(n146), .I3(n18277), .O(n839[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_16 (.CI(n18277), .I0(n840[13]), 
            .I1(n146), .CO(n767));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_15_lut (.I0(GND_net), .I1(n840[12]), 
            .I2(n141), .I3(n18276), .O(n839[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_15 (.CI(n18276), .I0(n840[12]), 
            .I1(n141), .CO(n18277));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_14_lut (.I0(GND_net), .I1(n840[11]), 
            .I2(n138_c), .I3(n18275), .O(n839[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_14 (.CI(n18275), .I0(n840[11]), 
            .I1(n138_c), .CO(n18276));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_13_lut (.I0(GND_net), .I1(n840[10]), 
            .I2(n135_c), .I3(n18274), .O(n839[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_13 (.CI(n18274), .I0(n840[10]), 
            .I1(n135_c), .CO(n18275));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_12_lut (.I0(GND_net), .I1(n840[9]), 
            .I2(n132_c), .I3(n18273), .O(n839[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_12 (.CI(n18273), .I0(n840[9]), 
            .I1(n132_c), .CO(n18274));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_11_lut (.I0(GND_net), .I1(n840[8]), 
            .I2(n129_c), .I3(n18272), .O(n839[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_11 (.CI(n18272), .I0(n840[8]), 
            .I1(n129_c), .CO(n18273));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_10_lut (.I0(GND_net), .I1(n840[7]), 
            .I2(n126_c), .I3(n18271), .O(n839[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_10 (.CI(n18271), .I0(n840[7]), 
            .I1(n126_c), .CO(n18272));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_9_lut (.I0(GND_net), .I1(n840[6]), 
            .I2(n123_c), .I3(n18270), .O(n839[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_9 (.CI(n18270), .I0(n840[6]), 
            .I1(n123_c), .CO(n18271));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_8_lut (.I0(GND_net), .I1(n840[5]), 
            .I2(n120_c), .I3(n18269), .O(n839[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_8 (.CI(n18269), .I0(n840[5]), 
            .I1(n120_c), .CO(n18270));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_7_lut (.I0(GND_net), .I1(n840[4]), 
            .I2(n117_c), .I3(n18268), .O(n839[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_7 (.CI(n18268), .I0(n840[4]), 
            .I1(n117_c), .CO(n18269));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_6_lut (.I0(GND_net), .I1(n840[3]), 
            .I2(n114_c), .I3(n18267), .O(n839[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_6 (.CI(n18267), .I0(n840[3]), 
            .I1(n114_c), .CO(n18268));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_5_lut (.I0(GND_net), .I1(n840[2]), 
            .I2(n111_c), .I3(n18266), .O(n839[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_5 (.CI(n18266), .I0(n840[2]), 
            .I1(n111_c), .CO(n18267));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_4_lut (.I0(GND_net), .I1(n840[1]), 
            .I2(n108_c), .I3(n18265), .O(n839[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_4 (.CI(n18265), .I0(n840[1]), 
            .I1(n108_c), .CO(n18266));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_3_lut (.I0(GND_net), .I1(n840[0]), 
            .I2(n105_c), .I3(n18264), .O(n839[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_3 (.CI(n18264), .I0(n840[0]), 
            .I1(n105_c), .CO(n18265));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n839[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18264));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_16_lut (.I0(GND_net), .I1(n839[13]), 
            .I2(n146), .I3(n18262), .O(n838[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_16 (.CI(n18262), .I0(n839[13]), 
            .I1(n146), .CO(n763));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_15_lut (.I0(GND_net), .I1(n839[12]), 
            .I2(n141), .I3(n18261), .O(n838[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_15 (.CI(n18261), .I0(n839[12]), 
            .I1(n141), .CO(n18262));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_14_lut (.I0(GND_net), .I1(n839[11]), 
            .I2(n138_c), .I3(n18260), .O(n838[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_14 (.CI(n18260), .I0(n839[11]), 
            .I1(n138_c), .CO(n18261));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_13_lut (.I0(GND_net), .I1(n839[10]), 
            .I2(n135_c), .I3(n18259), .O(n838[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_13 (.CI(n18259), .I0(n839[10]), 
            .I1(n135_c), .CO(n18260));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_12_lut (.I0(GND_net), .I1(n839[9]), 
            .I2(n132_c), .I3(n18258), .O(n838[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_12 (.CI(n18258), .I0(n839[9]), 
            .I1(n132_c), .CO(n18259));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_11_lut (.I0(GND_net), .I1(n839[8]), 
            .I2(n129_c), .I3(n18257), .O(n838[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_11 (.CI(n18257), .I0(n839[8]), 
            .I1(n129_c), .CO(n18258));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_10_lut (.I0(GND_net), .I1(n839[7]), 
            .I2(n126_c), .I3(n18256), .O(n838[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_10 (.CI(n18256), .I0(n839[7]), 
            .I1(n126_c), .CO(n18257));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_9_lut (.I0(GND_net), .I1(n839[6]), 
            .I2(n123_c), .I3(n18255), .O(n838[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_9 (.CI(n18255), .I0(n839[6]), 
            .I1(n123_c), .CO(n18256));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_8_lut (.I0(GND_net), .I1(n839[5]), 
            .I2(n120_c), .I3(n18254), .O(n838[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_8 (.CI(n18254), .I0(n839[5]), 
            .I1(n120_c), .CO(n18255));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_7_lut (.I0(GND_net), .I1(n839[4]), 
            .I2(n117_c), .I3(n18253), .O(n838[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_7 (.CI(n18253), .I0(n839[4]), 
            .I1(n117_c), .CO(n18254));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_6_lut (.I0(GND_net), .I1(n839[3]), 
            .I2(n114_c), .I3(n18252), .O(n838[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_6 (.CI(n18252), .I0(n839[3]), 
            .I1(n114_c), .CO(n18253));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_5_lut (.I0(GND_net), .I1(n839[2]), 
            .I2(n111_c), .I3(n18251), .O(n838[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_5 (.CI(n18251), .I0(n839[2]), 
            .I1(n111_c), .CO(n18252));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_4_lut (.I0(GND_net), .I1(n839[1]), 
            .I2(n108_c), .I3(n18250), .O(n838[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_4 (.CI(n18250), .I0(n839[1]), 
            .I1(n108_c), .CO(n18251));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_3_lut (.I0(GND_net), .I1(n839[0]), 
            .I2(n105_c), .I3(n18249), .O(n838[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_3 (.CI(n18249), .I0(n839[0]), 
            .I1(n105_c), .CO(n18250));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n838[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18249));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_16_lut (.I0(GND_net), .I1(n838[13]), 
            .I2(n146), .I3(n18247), .O(n837[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_16 (.CI(n18247), .I0(n838[13]), 
            .I1(n146), .CO(n759));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_15_lut (.I0(GND_net), .I1(n838[12]), 
            .I2(n141), .I3(n18246), .O(n837[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_15 (.CI(n18246), .I0(n838[12]), 
            .I1(n141), .CO(n18247));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_14_lut (.I0(GND_net), .I1(n838[11]), 
            .I2(n138_c), .I3(n18245), .O(n837[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_14 (.CI(n18245), .I0(n838[11]), 
            .I1(n138_c), .CO(n18246));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_13_lut (.I0(GND_net), .I1(n838[10]), 
            .I2(n135_c), .I3(n18244), .O(n837[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_13 (.CI(n18244), .I0(n838[10]), 
            .I1(n135_c), .CO(n18245));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_12_lut (.I0(GND_net), .I1(n838[9]), 
            .I2(n132_c), .I3(n18243), .O(n837[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_12 (.CI(n18243), .I0(n838[9]), 
            .I1(n132_c), .CO(n18244));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_11_lut (.I0(GND_net), .I1(n838[8]), 
            .I2(n129_c), .I3(n18242), .O(n837[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_11 (.CI(n18242), .I0(n838[8]), 
            .I1(n129_c), .CO(n18243));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_10_lut (.I0(GND_net), .I1(n838[7]), 
            .I2(n126_c), .I3(n18241), .O(n837[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_10 (.CI(n18241), .I0(n838[7]), 
            .I1(n126_c), .CO(n18242));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_9_lut (.I0(GND_net), .I1(n838[6]), 
            .I2(n123_c), .I3(n18240), .O(n837[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_9 (.CI(n18240), .I0(n838[6]), 
            .I1(n123_c), .CO(n18241));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_8_lut (.I0(GND_net), .I1(n838[5]), 
            .I2(n120_c), .I3(n18239), .O(n837[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_8 (.CI(n18239), .I0(n838[5]), 
            .I1(n120_c), .CO(n18240));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_7_lut (.I0(GND_net), .I1(n838[4]), 
            .I2(n117_c), .I3(n18238), .O(n837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_7 (.CI(n18238), .I0(n838[4]), 
            .I1(n117_c), .CO(n18239));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_6_lut (.I0(GND_net), .I1(n838[3]), 
            .I2(n114_c), .I3(n18237), .O(n837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_6 (.CI(n18237), .I0(n838[3]), 
            .I1(n114_c), .CO(n18238));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_5_lut (.I0(GND_net), .I1(n838[2]), 
            .I2(n111_c), .I3(n18236), .O(n837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_5 (.CI(n18236), .I0(n838[2]), 
            .I1(n111_c), .CO(n18237));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_4_lut (.I0(GND_net), .I1(n838[1]), 
            .I2(n108_c), .I3(n18235), .O(n837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_4 (.CI(n18235), .I0(n838[1]), 
            .I1(n108_c), .CO(n18236));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_3_lut (.I0(GND_net), .I1(n838[0]), 
            .I2(n105_c), .I3(n18234), .O(n837[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_3 (.CI(n18234), .I0(n838[0]), 
            .I1(n105_c), .CO(n18235));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n837[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18234));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_16_lut (.I0(GND_net), .I1(n837[13]), 
            .I2(n146), .I3(n18232), .O(n836[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_16 (.CI(n18232), .I0(n837[13]), 
            .I1(n146), .CO(n755));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_15_lut (.I0(GND_net), .I1(n837[12]), 
            .I2(n141), .I3(n18231), .O(n836[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_15 (.CI(n18231), .I0(n837[12]), 
            .I1(n141), .CO(n18232));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_14_lut (.I0(GND_net), .I1(n837[11]), 
            .I2(n138_c), .I3(n18230), .O(n836[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_14 (.CI(n18230), .I0(n837[11]), 
            .I1(n138_c), .CO(n18231));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_13_lut (.I0(GND_net), .I1(n837[10]), 
            .I2(n135_c), .I3(n18229), .O(n836[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_13 (.CI(n18229), .I0(n837[10]), 
            .I1(n135_c), .CO(n18230));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_12_lut (.I0(GND_net), .I1(n837[9]), 
            .I2(n132_c), .I3(n18228), .O(n836[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_12 (.CI(n18228), .I0(n837[9]), 
            .I1(n132_c), .CO(n18229));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_11_lut (.I0(GND_net), .I1(n837[8]), 
            .I2(n129_c), .I3(n18227), .O(n836[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_11 (.CI(n18227), .I0(n837[8]), 
            .I1(n129_c), .CO(n18228));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_10_lut (.I0(GND_net), .I1(n837[7]), 
            .I2(n126_c), .I3(n18226), .O(n836[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_10 (.CI(n18226), .I0(n837[7]), 
            .I1(n126_c), .CO(n18227));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_9_lut (.I0(GND_net), .I1(n837[6]), 
            .I2(n123_c), .I3(n18225), .O(n836[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_9 (.CI(n18225), .I0(n837[6]), 
            .I1(n123_c), .CO(n18226));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_8_lut (.I0(GND_net), .I1(n837[5]), 
            .I2(n120_c), .I3(n18224), .O(n836[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_8 (.CI(n18224), .I0(n837[5]), 
            .I1(n120_c), .CO(n18225));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n837[4]), 
            .I2(n117_c), .I3(n18223), .O(n836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_7 (.CI(n18223), .I0(n837[4]), 
            .I1(n117_c), .CO(n18224));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n837[3]), 
            .I2(n114_c), .I3(n18222), .O(n836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_6 (.CI(n18222), .I0(n837[3]), 
            .I1(n114_c), .CO(n18223));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n837[2]), 
            .I2(n111_c), .I3(n18221), .O(n836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_5 (.CI(n18221), .I0(n837[2]), 
            .I1(n111_c), .CO(n18222));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n837[1]), 
            .I2(n108_c), .I3(n18220), .O(n836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_4 (.CI(n18220), .I0(n837[1]), 
            .I1(n108_c), .CO(n18221));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n837[0]), 
            .I2(n105_c), .I3(n18219), .O(n836[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_3 (.CI(n18219), .I0(n837[0]), 
            .I1(n105_c), .CO(n18220));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n836[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18219));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_16_lut (.I0(GND_net), .I1(n836[13]), 
            .I2(n146), .I3(n18217), .O(n835[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_16 (.CI(n18217), .I0(n836[13]), 
            .I1(n146), .CO(n751));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_15_lut (.I0(GND_net), .I1(n836[12]), 
            .I2(n141), .I3(n18216), .O(n835[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_15 (.CI(n18216), .I0(n836[12]), 
            .I1(n141), .CO(n18217));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_14_lut (.I0(GND_net), .I1(n836[11]), 
            .I2(n138_c), .I3(n18215), .O(n835[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_14 (.CI(n18215), .I0(n836[11]), 
            .I1(n138_c), .CO(n18216));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_13_lut (.I0(GND_net), .I1(n836[10]), 
            .I2(n135_c), .I3(n18214), .O(n835[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_13 (.CI(n18214), .I0(n836[10]), 
            .I1(n135_c), .CO(n18215));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_12_lut (.I0(GND_net), .I1(n836[9]), 
            .I2(n132_c), .I3(n18213), .O(n835[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_12 (.CI(n18213), .I0(n836[9]), 
            .I1(n132_c), .CO(n18214));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_11_lut (.I0(GND_net), .I1(n836[8]), 
            .I2(n129_c), .I3(n18212), .O(n835[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_11 (.CI(n18212), .I0(n836[8]), 
            .I1(n129_c), .CO(n18213));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_10_lut (.I0(GND_net), .I1(n836[7]), 
            .I2(n126_c), .I3(n18211), .O(n835[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_10 (.CI(n18211), .I0(n836[7]), 
            .I1(n126_c), .CO(n18212));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_9_lut (.I0(GND_net), .I1(n836[6]), 
            .I2(n123_c), .I3(n18210), .O(n835[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_9 (.CI(n18210), .I0(n836[6]), 
            .I1(n123_c), .CO(n18211));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_8_lut (.I0(GND_net), .I1(n836[5]), 
            .I2(n120_c), .I3(n18209), .O(n835[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_8 (.CI(n18209), .I0(n836[5]), 
            .I1(n120_c), .CO(n18210));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_7_lut (.I0(GND_net), .I1(n836[4]), 
            .I2(n117_c), .I3(n18208), .O(n835[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_7 (.CI(n18208), .I0(n836[4]), 
            .I1(n117_c), .CO(n18209));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_6_lut (.I0(GND_net), .I1(n836[3]), 
            .I2(n114_c), .I3(n18207), .O(n835[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_6 (.CI(n18207), .I0(n836[3]), 
            .I1(n114_c), .CO(n18208));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_5_lut (.I0(GND_net), .I1(n836[2]), 
            .I2(n111_c), .I3(n18206), .O(n835[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_5 (.CI(n18206), .I0(n836[2]), 
            .I1(n111_c), .CO(n18207));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_4_lut (.I0(GND_net), .I1(n836[1]), 
            .I2(n108_c), .I3(n18205), .O(n835[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_4 (.CI(n18205), .I0(n836[1]), 
            .I1(n108_c), .CO(n18206));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_3_lut (.I0(GND_net), .I1(n836[0]), 
            .I2(n105_c), .I3(n18204), .O(n835[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_3 (.CI(n18204), .I0(n836[0]), 
            .I1(n105_c), .CO(n18205));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n835[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18204));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_16_lut (.I0(GND_net), .I1(n835[13]), 
            .I2(n146), .I3(n18202), .O(n834[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_16 (.CI(n18202), .I0(n835[13]), 
            .I1(n146), .CO(n747));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_15_lut (.I0(GND_net), .I1(n835[12]), 
            .I2(n141), .I3(n18201), .O(n834[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_15 (.CI(n18201), .I0(n835[12]), 
            .I1(n141), .CO(n18202));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_14_lut (.I0(GND_net), .I1(n835[11]), 
            .I2(n138_c), .I3(n18200), .O(n834[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_14 (.CI(n18200), .I0(n835[11]), 
            .I1(n138_c), .CO(n18201));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_13_lut (.I0(GND_net), .I1(n835[10]), 
            .I2(n135_c), .I3(n18199), .O(n834[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_13 (.CI(n18199), .I0(n835[10]), 
            .I1(n135_c), .CO(n18200));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_12_lut (.I0(GND_net), .I1(n835[9]), 
            .I2(n132_c), .I3(n18198), .O(n834[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_12 (.CI(n18198), .I0(n835[9]), 
            .I1(n132_c), .CO(n18199));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_11_lut (.I0(GND_net), .I1(n835[8]), 
            .I2(n129_c), .I3(n18197), .O(n834[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_11 (.CI(n18197), .I0(n835[8]), 
            .I1(n129_c), .CO(n18198));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_10_lut (.I0(GND_net), .I1(n835[7]), 
            .I2(n126_c), .I3(n18196), .O(n834[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_10 (.CI(n18196), .I0(n835[7]), 
            .I1(n126_c), .CO(n18197));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_9_lut (.I0(GND_net), .I1(n835[6]), 
            .I2(n123_c), .I3(n18195), .O(n834[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_9 (.CI(n18195), .I0(n835[6]), 
            .I1(n123_c), .CO(n18196));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_8_lut (.I0(GND_net), .I1(n835[5]), 
            .I2(n120_c), .I3(n18194), .O(n834[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_8 (.CI(n18194), .I0(n835[5]), 
            .I1(n120_c), .CO(n18195));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_7_lut (.I0(GND_net), .I1(n835[4]), 
            .I2(n117_c), .I3(n18193), .O(n834[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_7 (.CI(n18193), .I0(n835[4]), 
            .I1(n117_c), .CO(n18194));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_6_lut (.I0(GND_net), .I1(n835[3]), 
            .I2(n114_c), .I3(n18192), .O(n834[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_6 (.CI(n18192), .I0(n835[3]), 
            .I1(n114_c), .CO(n18193));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_5_lut (.I0(GND_net), .I1(n835[2]), 
            .I2(n111_c), .I3(n18191), .O(n834[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_5 (.CI(n18191), .I0(n835[2]), 
            .I1(n111_c), .CO(n18192));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_4_lut (.I0(GND_net), .I1(n835[1]), 
            .I2(n108_c), .I3(n18190), .O(n834[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_4 (.CI(n18190), .I0(n835[1]), 
            .I1(n108_c), .CO(n18191));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_3_lut (.I0(GND_net), .I1(n835[0]), 
            .I2(n105_c), .I3(n18189), .O(n834[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_3 (.CI(n18189), .I0(n835[0]), 
            .I1(n105_c), .CO(n18190));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n834[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18189));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_16_lut (.I0(GND_net), .I1(n834[13]), 
            .I2(n146), .I3(n18187), .O(n833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_16 (.CI(n18187), .I0(n834[13]), 
            .I1(n146), .CO(n743));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_15_lut (.I0(GND_net), .I1(n834[12]), 
            .I2(n141), .I3(n18186), .O(n833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_15 (.CI(n18186), .I0(n834[12]), 
            .I1(n141), .CO(n18187));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_14_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[11]), .I2(n138_c), .I3(n18185), .O(Switch_out1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_14 (.CI(n18185), .I0(n834[11]), 
            .I1(n138_c), .CO(n18186));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_13_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[10]), .I2(n135_c), .I3(n18184), .O(Switch_out1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_13 (.CI(n18184), .I0(n834[10]), 
            .I1(n135_c), .CO(n18185));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_12_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[9]), .I2(n132_c), .I3(n18183), .O(Switch_out1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_12 (.CI(n18183), .I0(n834[9]), 
            .I1(n132_c), .CO(n18184));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_11_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[8]), .I2(n129_c), .I3(n18182), .O(Switch_out1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_11 (.CI(n18182), .I0(n834[8]), 
            .I1(n129_c), .CO(n18183));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_10_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[7]), .I2(n126_c), .I3(n18181), .O(Switch_out1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_10 (.CI(n18181), .I0(n834[7]), 
            .I1(n126_c), .CO(n18182));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_9_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[6]), .I2(n123_c), .I3(n18180), .O(Switch_out1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_9 (.CI(n18180), .I0(n834[6]), 
            .I1(n123_c), .CO(n18181));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_8_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[5]), .I2(n120_c), .I3(n18179), .O(Switch_out1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_8 (.CI(n18179), .I0(n834[5]), 
            .I1(n120_c), .CO(n18180));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_7_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[4]), .I2(n117_c), .I3(n18178), .O(Switch_out1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_7 (.CI(n18178), .I0(n834[4]), 
            .I1(n117_c), .CO(n18179));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_6_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[3]), .I2(n114_c), .I3(n18177), .O(Switch_out1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_6 (.CI(n18177), .I0(n834[3]), 
            .I1(n114_c), .CO(n18178));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_5_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[2]), .I2(n111_c), .I3(n18176), .O(Switch_out1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_5 (.CI(n18176), .I0(n834[2]), 
            .I1(n111_c), .CO(n18177));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_4_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[1]), .I2(n108_c), .I3(n18175), .O(Switch_out1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_4 (.CI(n18175), .I0(n834[1]), 
            .I1(n108_c), .CO(n18176));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_3_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834[0]), .I2(n105_c), .I3(n18174), .O(Switch_out1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_3 (.CI(n18174), .I0(n834[0]), 
            .I1(n105_c), .CO(n18175));
    SB_CARRY Error_sub_temp_31__I_0_add_562_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n18174));
    SB_LUT4 add_4259_17_lut (.I0(Not_Equal_relop1_N_201), .I1(n796), .I2(n795), 
            .I3(n18159), .O(Switch_out1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4259_16_lut (.I0(Not_Equal_relop1_N_201), .I1(n846[14]), 
            .I2(n791), .I3(n18158), .O(Switch_out1[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_16 (.CI(n18158), .I0(n846[14]), .I1(n791), .CO(n18159));
    SB_LUT4 add_4259_15_lut (.I0(Not_Equal_relop1_N_201), .I1(n845[14]), 
            .I2(n787), .I3(n18157), .O(Switch_out1[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_15 (.CI(n18157), .I0(n845[14]), .I1(n787), .CO(n18158));
    SB_LUT4 add_4259_14_lut (.I0(Not_Equal_relop1_N_201), .I1(n844[14]), 
            .I2(n783), .I3(n18156), .O(Switch_out1[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_14 (.CI(n18156), .I0(n844[14]), .I1(n783), .CO(n18157));
    SB_LUT4 add_4259_13_lut (.I0(Not_Equal_relop1_N_201), .I1(n843[14]), 
            .I2(n779), .I3(n18155), .O(Switch_out1[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_13 (.CI(n18155), .I0(n843[14]), .I1(n779), .CO(n18156));
    SB_LUT4 add_4259_12_lut (.I0(Not_Equal_relop1_N_201), .I1(n842_adj_806[14]), 
            .I2(n775_adj_590), .I3(n18154), .O(Switch_out1[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_12 (.CI(n18154), .I0(n842_adj_806[14]), .I1(n775_adj_590), 
            .CO(n18155));
    SB_LUT4 add_4259_11_lut (.I0(Not_Equal_relop1_N_201), .I1(n841_adj_807[14]), 
            .I2(n771), .I3(n18153), .O(Switch_out1[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_11 (.CI(n18153), .I0(n841_adj_807[14]), .I1(n771), 
            .CO(n18154));
    SB_LUT4 add_4259_10_lut (.I0(Not_Equal_relop1_N_201), .I1(n840[14]), 
            .I2(n767), .I3(n18152), .O(Switch_out1[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_10 (.CI(n18152), .I0(n840[14]), .I1(n767), .CO(n18153));
    SB_LUT4 add_4259_9_lut (.I0(Not_Equal_relop1_N_201), .I1(n839[14]), 
            .I2(n763), .I3(n18151), .O(Switch_out1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_9 (.CI(n18151), .I0(n839[14]), .I1(n763), .CO(n18152));
    SB_LUT4 add_4259_8_lut (.I0(Not_Equal_relop1_N_201), .I1(n838[14]), 
            .I2(n759), .I3(n18150), .O(Switch_out1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_8 (.CI(n18150), .I0(n838[14]), .I1(n759), .CO(n18151));
    SB_LUT4 add_4259_7_lut (.I0(Not_Equal_relop1_N_201), .I1(n837[14]), 
            .I2(n755), .I3(n18149), .O(Switch_out1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4259_6_lut (.I0(Not_Equal_relop1_N_201), .I1(n836[14]), 
            .I2(n751), .I3(n18148), .O(Switch_out1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_6 (.CI(n18148), .I0(n836[14]), .I1(n751), .CO(n18149));
    SB_CARRY add_4259_7 (.CI(n18149), .I0(n837[14]), .I1(n755), .CO(n18150));
    SB_LUT4 add_4259_5_lut (.I0(Not_Equal_relop1_N_201), .I1(n835[14]), 
            .I2(n747), .I3(n18147), .O(Switch_out1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_5 (.CI(n18147), .I0(n835[14]), .I1(n747), .CO(n18148));
    SB_LUT4 add_4259_4_lut (.I0(Not_Equal_relop1_N_201), .I1(n834[14]), 
            .I2(n743), .I3(n18146), .O(Switch_out1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_4 (.CI(n18146), .I0(n834[14]), .I1(n743), .CO(n18147));
    SB_LUT4 add_4259_3_lut (.I0(Not_Equal_relop1_N_201), .I1(n833[14]), 
            .I2(n8356), .I3(n18145), .O(Switch_out1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_3 (.CI(n18145), .I0(n833[14]), .I1(n8356), .CO(n18146));
    SB_LUT4 add_4259_2_lut (.I0(Not_Equal_relop1_N_201), .I1(\Error_sub_temp[31] ), 
            .I2(\Product_mul_temp[26] ), .I3(n18144), .O(Switch_out1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4259_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4259_2 (.CI(n18144), .I0(\Error_sub_temp[31] ), .I1(\Product_mul_temp[26] ), 
            .CO(n18145));
    SB_CARRY add_4259_1 (.CI(GND_net), .I0(n832[14]), .I1(n832[14]), .CO(n18144));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_16_lut (.I0(GND_net), .I1(n841[11]), 
            .I2(n769_c), .I3(n18120), .O(n840_adj_808[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_16 (.CI(n18120), .I0(n841[11]), 
            .I1(n769_c), .CO(n771_adj_598));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_15_lut (.I0(GND_net), .I1(n841[11]), 
            .I2(n123_c), .I3(n18119), .O(n840_adj_808[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_15 (.CI(n18119), .I0(n841[11]), 
            .I1(n123_c), .CO(n18120));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_14_lut (.I0(GND_net), .I1(n841[11]), 
            .I2(n123_c), .I3(n18118), .O(n840_adj_808[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_14 (.CI(n18118), .I0(n841[11]), 
            .I1(n123_c), .CO(n18119));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_13_lut (.I0(GND_net), .I1(n841[10]), 
            .I2(n123_c), .I3(n18117), .O(n840_adj_808[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_13 (.CI(n18117), .I0(n841[10]), 
            .I1(n123_c), .CO(n18118));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_12_lut (.I0(GND_net), .I1(n841[9]), 
            .I2(n123_c), .I3(n18116), .O(n840_adj_808[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_12 (.CI(n18116), .I0(n841[9]), 
            .I1(n123_c), .CO(n18117));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_11_lut (.I0(GND_net), .I1(n841[8]), 
            .I2(n123_c), .I3(n18115), .O(n840_adj_808[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_11 (.CI(n18115), .I0(n841[8]), 
            .I1(n123_c), .CO(n18116));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_10_lut (.I0(GND_net), .I1(n841[7]), 
            .I2(n123_c), .I3(n18114), .O(n840_adj_808[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_10 (.CI(n18114), .I0(n841[7]), 
            .I1(n123_c), .CO(n18115));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_9_lut (.I0(GND_net), .I1(n841[6]), 
            .I2(n123_c), .I3(n18113), .O(n840_adj_808[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_9 (.CI(n18113), .I0(n841[6]), 
            .I1(n123_c), .CO(n18114));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_8_lut (.I0(GND_net), .I1(n841[5]), 
            .I2(n123_c), .I3(n18112), .O(n840_adj_808[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_8 (.CI(n18112), .I0(n841[5]), 
            .I1(n123_c), .CO(n18113));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_7_lut (.I0(GND_net), .I1(n841[4]), 
            .I2(n123_c), .I3(n18111), .O(n840_adj_808[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_7 (.CI(n18111), .I0(n841[4]), 
            .I1(n123_c), .CO(n18112));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_6_lut (.I0(GND_net), .I1(n841[3]), 
            .I2(n123_c), .I3(n18110), .O(n840_adj_808[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_6 (.CI(n18110), .I0(n841[3]), 
            .I1(n123_c), .CO(n18111));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_5_lut (.I0(GND_net), .I1(n841[2]), 
            .I2(n123_c), .I3(n18109), .O(n840_adj_808[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_5 (.CI(n18109), .I0(n841[2]), 
            .I1(n123_c), .CO(n18110));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_4_lut (.I0(GND_net), .I1(n841[1]), 
            .I2(n123_c), .I3(n18108), .O(n840_adj_808[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_4 (.CI(n18108), .I0(n841[1]), 
            .I1(n123_c), .CO(n18109));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_3_lut (.I0(GND_net), .I1(n841[0]), 
            .I2(n123_c), .I3(n18107), .O(n840_adj_808[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_3 (.CI(n18107), .I0(n841[0]), 
            .I1(n123_c), .CO(n18108));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_2_lut (.I0(GND_net), .I1(n126_c), 
            .I2(n123_c), .I3(GND_net), .O(n840_adj_808[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_2 (.CI(GND_net), .I0(n126_c), 
            .I1(n123_c), .CO(n18107));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_16_lut (.I0(GND_net), .I1(n840_adj_808[13]), 
            .I2(n765_c), .I3(n18105), .O(n839_adj_809[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_16 (.CI(n18105), .I0(n840_adj_808[13]), 
            .I1(n765_c), .CO(n767_adj_620));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_15_lut (.I0(GND_net), .I1(n840_adj_808[12]), 
            .I2(n120_c), .I3(n18104), .O(n839_adj_809[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_15 (.CI(n18104), .I0(n840_adj_808[12]), 
            .I1(n120_c), .CO(n18105));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_14_lut (.I0(GND_net), .I1(n840_adj_808[11]), 
            .I2(n120_c), .I3(n18103), .O(n839_adj_809[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_14 (.CI(n18103), .I0(n840_adj_808[11]), 
            .I1(n120_c), .CO(n18104));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_13_lut (.I0(GND_net), .I1(n840_adj_808[10]), 
            .I2(n120_c), .I3(n18102), .O(n839_adj_809[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_13 (.CI(n18102), .I0(n840_adj_808[10]), 
            .I1(n120_c), .CO(n18103));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_12_lut (.I0(GND_net), .I1(n840_adj_808[9]), 
            .I2(n120_c), .I3(n18101), .O(n839_adj_809[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_12 (.CI(n18101), .I0(n840_adj_808[9]), 
            .I1(n120_c), .CO(n18102));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_11_lut (.I0(GND_net), .I1(n840_adj_808[8]), 
            .I2(n120_c), .I3(n18100), .O(n839_adj_809[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_11 (.CI(n18100), .I0(n840_adj_808[8]), 
            .I1(n120_c), .CO(n18101));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_10_lut (.I0(GND_net), .I1(n840_adj_808[7]), 
            .I2(n120_c), .I3(n18099), .O(n839_adj_809[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_10 (.CI(n18099), .I0(n840_adj_808[7]), 
            .I1(n120_c), .CO(n18100));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_9_lut (.I0(GND_net), .I1(n840_adj_808[6]), 
            .I2(n120_c), .I3(n18098), .O(n839_adj_809[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_9 (.CI(n18098), .I0(n840_adj_808[6]), 
            .I1(n120_c), .CO(n18099));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_8_lut (.I0(GND_net), .I1(n840_adj_808[5]), 
            .I2(n120_c), .I3(n18097), .O(n839_adj_809[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_8 (.CI(n18097), .I0(n840_adj_808[5]), 
            .I1(n120_c), .CO(n18098));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_7_lut (.I0(GND_net), .I1(n840_adj_808[4]), 
            .I2(n120_c), .I3(n18096), .O(n839_adj_809[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_7 (.CI(n18096), .I0(n840_adj_808[4]), 
            .I1(n120_c), .CO(n18097));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_6_lut (.I0(GND_net), .I1(n840_adj_808[3]), 
            .I2(n120_c), .I3(n18095), .O(n839_adj_809[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_6 (.CI(n18095), .I0(n840_adj_808[3]), 
            .I1(n120_c), .CO(n18096));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_5_lut (.I0(GND_net), .I1(n840_adj_808[2]), 
            .I2(n120_c), .I3(n18094), .O(n839_adj_809[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_5 (.CI(n18094), .I0(n840_adj_808[2]), 
            .I1(n120_c), .CO(n18095));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_4_lut (.I0(GND_net), .I1(n840_adj_808[1]), 
            .I2(n120_c), .I3(n18093), .O(n839_adj_809[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_4 (.CI(n18093), .I0(n840_adj_808[1]), 
            .I1(n120_c), .CO(n18094));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_3_lut (.I0(GND_net), .I1(n840_adj_808[0]), 
            .I2(n120_c), .I3(n18092), .O(n839_adj_809[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_3 (.CI(n18092), .I0(n840_adj_808[0]), 
            .I1(n120_c), .CO(n18093));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_2_lut (.I0(GND_net), .I1(n123_c), 
            .I2(n120_c), .I3(GND_net), .O(n839_adj_809[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_2 (.CI(GND_net), .I0(n123_c), 
            .I1(n120_c), .CO(n18092));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_16_lut (.I0(GND_net), .I1(n839_adj_809[13]), 
            .I2(n761_c), .I3(n18090), .O(n838_adj_810[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_16 (.CI(n18090), .I0(n839_adj_809[13]), 
            .I1(n761_c), .CO(n763_adj_636));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_15_lut (.I0(GND_net), .I1(n839_adj_809[12]), 
            .I2(n117_c), .I3(n18089), .O(n838_adj_810[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_15 (.CI(n18089), .I0(n839_adj_809[12]), 
            .I1(n117_c), .CO(n18090));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_14_lut (.I0(GND_net), .I1(n839_adj_809[11]), 
            .I2(n117_c), .I3(n18088), .O(n838_adj_810[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_14 (.CI(n18088), .I0(n839_adj_809[11]), 
            .I1(n117_c), .CO(n18089));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_13_lut (.I0(GND_net), .I1(n839_adj_809[10]), 
            .I2(n117_c), .I3(n18087), .O(n838_adj_810[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_13 (.CI(n18087), .I0(n839_adj_809[10]), 
            .I1(n117_c), .CO(n18088));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_12_lut (.I0(GND_net), .I1(n839_adj_809[9]), 
            .I2(n117_c), .I3(n18086), .O(n838_adj_810[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_12 (.CI(n18086), .I0(n839_adj_809[9]), 
            .I1(n117_c), .CO(n18087));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_11_lut (.I0(GND_net), .I1(n839_adj_809[8]), 
            .I2(n117_c), .I3(n18085), .O(n838_adj_810[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_11 (.CI(n18085), .I0(n839_adj_809[8]), 
            .I1(n117_c), .CO(n18086));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_10_lut (.I0(GND_net), .I1(n839_adj_809[7]), 
            .I2(n117_c), .I3(n18084), .O(n838_adj_810[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_10 (.CI(n18084), .I0(n839_adj_809[7]), 
            .I1(n117_c), .CO(n18085));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_9_lut (.I0(GND_net), .I1(n839_adj_809[6]), 
            .I2(n117_c), .I3(n18083), .O(n838_adj_810[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_9 (.CI(n18083), .I0(n839_adj_809[6]), 
            .I1(n117_c), .CO(n18084));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_8_lut (.I0(GND_net), .I1(n839_adj_809[5]), 
            .I2(n117_c), .I3(n18082), .O(n838_adj_810[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_8 (.CI(n18082), .I0(n839_adj_809[5]), 
            .I1(n117_c), .CO(n18083));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_7_lut (.I0(GND_net), .I1(n839_adj_809[4]), 
            .I2(n117_c), .I3(n18081), .O(n838_adj_810[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_7 (.CI(n18081), .I0(n839_adj_809[4]), 
            .I1(n117_c), .CO(n18082));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_6_lut (.I0(GND_net), .I1(n839_adj_809[3]), 
            .I2(n117_c), .I3(n18080), .O(n838_adj_810[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_6 (.CI(n18080), .I0(n839_adj_809[3]), 
            .I1(n117_c), .CO(n18081));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_5_lut (.I0(GND_net), .I1(n839_adj_809[2]), 
            .I2(n117_c), .I3(n18079), .O(n838_adj_810[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_5 (.CI(n18079), .I0(n839_adj_809[2]), 
            .I1(n117_c), .CO(n18080));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_4_lut (.I0(GND_net), .I1(n839_adj_809[1]), 
            .I2(n117_c), .I3(n18078), .O(n838_adj_810[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_4 (.CI(n18078), .I0(n839_adj_809[1]), 
            .I1(n117_c), .CO(n18079));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_3_lut (.I0(GND_net), .I1(n839_adj_809[0]), 
            .I2(n117_c), .I3(n18077), .O(n838_adj_810[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_3 (.CI(n18077), .I0(n839_adj_809[0]), 
            .I1(n117_c), .CO(n18078));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_2_lut (.I0(GND_net), .I1(n120_c), 
            .I2(n117_c), .I3(GND_net), .O(n838_adj_810[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_2 (.CI(GND_net), .I0(n120_c), 
            .I1(n117_c), .CO(n18077));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_16_lut (.I0(GND_net), .I1(n838_adj_810[13]), 
            .I2(n757_c), .I3(n18075), .O(n837_adj_811[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_16 (.CI(n18075), .I0(n838_adj_810[13]), 
            .I1(n757_c), .CO(n759_adj_652));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_15_lut (.I0(GND_net), .I1(n838_adj_810[12]), 
            .I2(n114_c), .I3(n18074), .O(n837_adj_811[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_15 (.CI(n18074), .I0(n838_adj_810[12]), 
            .I1(n114_c), .CO(n18075));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_14_lut (.I0(GND_net), .I1(n838_adj_810[11]), 
            .I2(n114_c), .I3(n18073), .O(n837_adj_811[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_14 (.CI(n18073), .I0(n838_adj_810[11]), 
            .I1(n114_c), .CO(n18074));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_13_lut (.I0(GND_net), .I1(n838_adj_810[10]), 
            .I2(n114_c), .I3(n18072), .O(n837_adj_811[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_13 (.CI(n18072), .I0(n838_adj_810[10]), 
            .I1(n114_c), .CO(n18073));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_12_lut (.I0(GND_net), .I1(n838_adj_810[9]), 
            .I2(n114_c), .I3(n18071), .O(n837_adj_811[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_12 (.CI(n18071), .I0(n838_adj_810[9]), 
            .I1(n114_c), .CO(n18072));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_11_lut (.I0(GND_net), .I1(n838_adj_810[8]), 
            .I2(n114_c), .I3(n18070), .O(n837_adj_811[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_11 (.CI(n18070), .I0(n838_adj_810[8]), 
            .I1(n114_c), .CO(n18071));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_10_lut (.I0(GND_net), .I1(n838_adj_810[7]), 
            .I2(n114_c), .I3(n18069), .O(n837_adj_811[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_10 (.CI(n18069), .I0(n838_adj_810[7]), 
            .I1(n114_c), .CO(n18070));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_9_lut (.I0(GND_net), .I1(n838_adj_810[6]), 
            .I2(n114_c), .I3(n18068), .O(n837_adj_811[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_9 (.CI(n18068), .I0(n838_adj_810[6]), 
            .I1(n114_c), .CO(n18069));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_8_lut (.I0(GND_net), .I1(n838_adj_810[5]), 
            .I2(n114_c), .I3(n18067), .O(n837_adj_811[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_8 (.CI(n18067), .I0(n838_adj_810[5]), 
            .I1(n114_c), .CO(n18068));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_7_lut (.I0(GND_net), .I1(n838_adj_810[4]), 
            .I2(n114_c), .I3(n18066), .O(n837_adj_811[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_7 (.CI(n18066), .I0(n838_adj_810[4]), 
            .I1(n114_c), .CO(n18067));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_6_lut (.I0(GND_net), .I1(n838_adj_810[3]), 
            .I2(n114_c), .I3(n18065), .O(n837_adj_811[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_6 (.CI(n18065), .I0(n838_adj_810[3]), 
            .I1(n114_c), .CO(n18066));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_5_lut (.I0(GND_net), .I1(n838_adj_810[2]), 
            .I2(n114_c), .I3(n18064), .O(n837_adj_811[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_5 (.CI(n18064), .I0(n838_adj_810[2]), 
            .I1(n114_c), .CO(n18065));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_4_lut (.I0(GND_net), .I1(n838_adj_810[1]), 
            .I2(n114_c), .I3(n18063), .O(n837_adj_811[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_4 (.CI(n18063), .I0(n838_adj_810[1]), 
            .I1(n114_c), .CO(n18064));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_3_lut (.I0(GND_net), .I1(n838_adj_810[0]), 
            .I2(n114_c), .I3(n18062), .O(n837_adj_811[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_3 (.CI(n18062), .I0(n838_adj_810[0]), 
            .I1(n114_c), .CO(n18063));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_2_lut (.I0(GND_net), .I1(n117_c), 
            .I2(n114_c), .I3(GND_net), .O(n837_adj_811[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_2 (.CI(GND_net), .I0(n117_c), 
            .I1(n114_c), .CO(n18062));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_16_lut (.I0(GND_net), .I1(n837_adj_811[13]), 
            .I2(n753_c), .I3(n18060), .O(n836_adj_812[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_16 (.CI(n18060), .I0(n837_adj_811[13]), 
            .I1(n753_c), .CO(n755_adj_668));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_15_lut (.I0(GND_net), .I1(n837_adj_811[12]), 
            .I2(n111_c), .I3(n18059), .O(n836_adj_812[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_15 (.CI(n18059), .I0(n837_adj_811[12]), 
            .I1(n111_c), .CO(n18060));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_14_lut (.I0(GND_net), .I1(n837_adj_811[11]), 
            .I2(n111_c), .I3(n18058), .O(n836_adj_812[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_14 (.CI(n18058), .I0(n837_adj_811[11]), 
            .I1(n111_c), .CO(n18059));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_13_lut (.I0(GND_net), .I1(n837_adj_811[10]), 
            .I2(n111_c), .I3(n18057), .O(n836_adj_812[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_13 (.CI(n18057), .I0(n837_adj_811[10]), 
            .I1(n111_c), .CO(n18058));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_12_lut (.I0(GND_net), .I1(n837_adj_811[9]), 
            .I2(n111_c), .I3(n18056), .O(n836_adj_812[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_12 (.CI(n18056), .I0(n837_adj_811[9]), 
            .I1(n111_c), .CO(n18057));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_11_lut (.I0(GND_net), .I1(n837_adj_811[8]), 
            .I2(n111_c), .I3(n18055), .O(n836_adj_812[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_11 (.CI(n18055), .I0(n837_adj_811[8]), 
            .I1(n111_c), .CO(n18056));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_10_lut (.I0(GND_net), .I1(n837_adj_811[7]), 
            .I2(n111_c), .I3(n18054), .O(n836_adj_812[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_10 (.CI(n18054), .I0(n837_adj_811[7]), 
            .I1(n111_c), .CO(n18055));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_9_lut (.I0(GND_net), .I1(n837_adj_811[6]), 
            .I2(n111_c), .I3(n18053), .O(n836_adj_812[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_9 (.CI(n18053), .I0(n837_adj_811[6]), 
            .I1(n111_c), .CO(n18054));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_8_lut (.I0(GND_net), .I1(n837_adj_811[5]), 
            .I2(n111_c), .I3(n18052), .O(n836_adj_812[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_8 (.CI(n18052), .I0(n837_adj_811[5]), 
            .I1(n111_c), .CO(n18053));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_7_lut (.I0(GND_net), .I1(n837_adj_811[4]), 
            .I2(n111_c), .I3(n18051), .O(n836_adj_812[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_7 (.CI(n18051), .I0(n837_adj_811[4]), 
            .I1(n111_c), .CO(n18052));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_6_lut (.I0(GND_net), .I1(n837_adj_811[3]), 
            .I2(n111_c), .I3(n18050), .O(n836_adj_812[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_6 (.CI(n18050), .I0(n837_adj_811[3]), 
            .I1(n111_c), .CO(n18051));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_5_lut (.I0(GND_net), .I1(n837_adj_811[2]), 
            .I2(n111_c), .I3(n18049), .O(n836_adj_812[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_5 (.CI(n18049), .I0(n837_adj_811[2]), 
            .I1(n111_c), .CO(n18050));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_4_lut (.I0(GND_net), .I1(n837_adj_811[1]), 
            .I2(n111_c), .I3(n18048), .O(n836_adj_812[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_4 (.CI(n18048), .I0(n837_adj_811[1]), 
            .I1(n111_c), .CO(n18049));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_3_lut (.I0(GND_net), .I1(n837_adj_811[0]), 
            .I2(n111_c), .I3(n18047), .O(n836_adj_812[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_3 (.CI(n18047), .I0(n837_adj_811[0]), 
            .I1(n111_c), .CO(n18048));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_2_lut (.I0(GND_net), .I1(n114_c), 
            .I2(n111_c), .I3(GND_net), .O(n836_adj_812[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_2 (.CI(GND_net), .I0(n114_c), 
            .I1(n111_c), .CO(n18047));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_16_lut (.I0(GND_net), .I1(n836_adj_812[13]), 
            .I2(n749_c), .I3(n18045), .O(n835_adj_813[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_16 (.CI(n18045), .I0(n836_adj_812[13]), 
            .I1(n749_c), .CO(n751_adj_684));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_15_lut (.I0(GND_net), .I1(n836_adj_812[12]), 
            .I2(n108_c), .I3(n18044), .O(n835_adj_813[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_15 (.CI(n18044), .I0(n836_adj_812[12]), 
            .I1(n108_c), .CO(n18045));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_14_lut (.I0(GND_net), .I1(n836_adj_812[11]), 
            .I2(n108_c), .I3(n18043), .O(n835_adj_813[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_14 (.CI(n18043), .I0(n836_adj_812[11]), 
            .I1(n108_c), .CO(n18044));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_13_lut (.I0(GND_net), .I1(n836_adj_812[10]), 
            .I2(n108_c), .I3(n18042), .O(n835_adj_813[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_13 (.CI(n18042), .I0(n836_adj_812[10]), 
            .I1(n108_c), .CO(n18043));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_12_lut (.I0(GND_net), .I1(n836_adj_812[9]), 
            .I2(n108_c), .I3(n18041), .O(n835_adj_813[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_12 (.CI(n18041), .I0(n836_adj_812[9]), 
            .I1(n108_c), .CO(n18042));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_11_lut (.I0(GND_net), .I1(n836_adj_812[8]), 
            .I2(n108_c), .I3(n18040), .O(n835_adj_813[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_11 (.CI(n18040), .I0(n836_adj_812[8]), 
            .I1(n108_c), .CO(n18041));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_10_lut (.I0(GND_net), .I1(n836_adj_812[7]), 
            .I2(n108_c), .I3(n18039), .O(n835_adj_813[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_10 (.CI(n18039), .I0(n836_adj_812[7]), 
            .I1(n108_c), .CO(n18040));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_9_lut (.I0(GND_net), .I1(n836_adj_812[6]), 
            .I2(n108_c), .I3(n18038), .O(n835_adj_813[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_9 (.CI(n18038), .I0(n836_adj_812[6]), 
            .I1(n108_c), .CO(n18039));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_8_lut (.I0(GND_net), .I1(n836_adj_812[5]), 
            .I2(n108_c), .I3(n18037), .O(n835_adj_813[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_8 (.CI(n18037), .I0(n836_adj_812[5]), 
            .I1(n108_c), .CO(n18038));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_7_lut (.I0(GND_net), .I1(n836_adj_812[4]), 
            .I2(n108_c), .I3(n18036), .O(n835_adj_813[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_7 (.CI(n18036), .I0(n836_adj_812[4]), 
            .I1(n108_c), .CO(n18037));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_6_lut (.I0(GND_net), .I1(n836_adj_812[3]), 
            .I2(n108_c), .I3(n18035), .O(n835_adj_813[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_6 (.CI(n18035), .I0(n836_adj_812[3]), 
            .I1(n108_c), .CO(n18036));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_5_lut (.I0(GND_net), .I1(n836_adj_812[2]), 
            .I2(n108_c), .I3(n18034), .O(n835_adj_813[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_5 (.CI(n18034), .I0(n836_adj_812[2]), 
            .I1(n108_c), .CO(n18035));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_4_lut (.I0(GND_net), .I1(n836_adj_812[1]), 
            .I2(n108_c), .I3(n18033), .O(n835_adj_813[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_4 (.CI(n18033), .I0(n836_adj_812[1]), 
            .I1(n108_c), .CO(n18034));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_3_lut (.I0(GND_net), .I1(n836_adj_812[0]), 
            .I2(n108_c), .I3(n18032), .O(n835_adj_813[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_3 (.CI(n18032), .I0(n836_adj_812[0]), 
            .I1(n108_c), .CO(n18033));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_2_lut (.I0(GND_net), .I1(n111_c), 
            .I2(n108_c), .I3(GND_net), .O(n835_adj_813[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_2 (.CI(GND_net), .I0(n111_c), 
            .I1(n108_c), .CO(n18032));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_16_lut (.I0(GND_net), .I1(n835_adj_813[13]), 
            .I2(n745_c), .I3(n18030), .O(n834_adj_814[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_16 (.CI(n18030), .I0(n835_adj_813[13]), 
            .I1(n745_c), .CO(n747_adj_700));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_15_lut (.I0(GND_net), .I1(n835_adj_813[12]), 
            .I2(n105_c), .I3(n18029), .O(n834_adj_814[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_15 (.CI(n18029), .I0(n835_adj_813[12]), 
            .I1(n105_c), .CO(n18030));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_14_lut (.I0(GND_net), .I1(n835_adj_813[11]), 
            .I2(n105_c), .I3(n18028), .O(n834_adj_814[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_14 (.CI(n18028), .I0(n835_adj_813[11]), 
            .I1(n105_c), .CO(n18029));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_13_lut (.I0(GND_net), .I1(n835_adj_813[10]), 
            .I2(n105_c), .I3(n18027), .O(n834_adj_814[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_13 (.CI(n18027), .I0(n835_adj_813[10]), 
            .I1(n105_c), .CO(n18028));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_12_lut (.I0(GND_net), .I1(n835_adj_813[9]), 
            .I2(n105_c), .I3(n18026), .O(n834_adj_814[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_12 (.CI(n18026), .I0(n835_adj_813[9]), 
            .I1(n105_c), .CO(n18027));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_11_lut (.I0(GND_net), .I1(n835_adj_813[8]), 
            .I2(n105_c), .I3(n18025), .O(n834_adj_814[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_11 (.CI(n18025), .I0(n835_adj_813[8]), 
            .I1(n105_c), .CO(n18026));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_10_lut (.I0(GND_net), .I1(n835_adj_813[7]), 
            .I2(n105_c), .I3(n18024), .O(n834_adj_814[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_10 (.CI(n18024), .I0(n835_adj_813[7]), 
            .I1(n105_c), .CO(n18025));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_9_lut (.I0(GND_net), .I1(n835_adj_813[6]), 
            .I2(n105_c), .I3(n18023), .O(n834_adj_814[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_9 (.CI(n18023), .I0(n835_adj_813[6]), 
            .I1(n105_c), .CO(n18024));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_8_lut (.I0(GND_net), .I1(n835_adj_813[5]), 
            .I2(n105_c), .I3(n18022), .O(n834_adj_814[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_8 (.CI(n18022), .I0(n835_adj_813[5]), 
            .I1(n105_c), .CO(n18023));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_7_lut (.I0(GND_net), .I1(n835_adj_813[4]), 
            .I2(n105_c), .I3(n18021), .O(n834_adj_814[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_7 (.CI(n18021), .I0(n835_adj_813[4]), 
            .I1(n105_c), .CO(n18022));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_6_lut (.I0(GND_net), .I1(n835_adj_813[3]), 
            .I2(n105_c), .I3(n18020), .O(n834_adj_814[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_6 (.CI(n18020), .I0(n835_adj_813[3]), 
            .I1(n105_c), .CO(n18021));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_5_lut (.I0(GND_net), .I1(n835_adj_813[2]), 
            .I2(n105_c), .I3(n18019), .O(n834_adj_814[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_5 (.CI(n18019), .I0(n835_adj_813[2]), 
            .I1(n105_c), .CO(n18020));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_4_lut (.I0(GND_net), .I1(n835_adj_813[1]), 
            .I2(n105_c), .I3(n18018), .O(n834_adj_814[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_4 (.CI(n18018), .I0(n835_adj_813[1]), 
            .I1(n105_c), .CO(n18019));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_3_lut (.I0(GND_net), .I1(n835_adj_813[0]), 
            .I2(n105_c), .I3(n18017), .O(n834_adj_814[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_3 (.CI(n18017), .I0(n835_adj_813[0]), 
            .I1(n105_c), .CO(n18018));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_2_lut (.I0(GND_net), .I1(n108_c), 
            .I2(n105_c), .I3(GND_net), .O(n834_adj_814[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_2 (.CI(GND_net), .I0(n108_c), 
            .I1(n105_c), .CO(n18017));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_16_lut (.I0(GND_net), .I1(n834_adj_814[13]), 
            .I2(n741_c), .I3(n18015), .O(n833_adj_815[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_16 (.CI(n18015), .I0(n834_adj_814[13]), 
            .I1(n741_c), .CO(n743_adj_716));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_15_lut (.I0(GND_net), .I1(n834_adj_814[12]), 
            .I2(n102_c), .I3(n18014), .O(n833_adj_815[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_15 (.CI(n18014), .I0(n834_adj_814[12]), 
            .I1(n102_c), .CO(n18015));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_14_lut (.I0(GND_net), .I1(n834_adj_814[11]), 
            .I2(n102_c), .I3(n18013), .O(n833_adj_815[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_14 (.CI(n18013), .I0(n834_adj_814[11]), 
            .I1(n102_c), .CO(n18014));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_13_lut (.I0(GND_net), .I1(n834_adj_814[10]), 
            .I2(n102_c), .I3(n18012), .O(n833_adj_815[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_13 (.CI(n18012), .I0(n834_adj_814[10]), 
            .I1(n102_c), .CO(n18013));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_12_lut (.I0(GND_net), .I1(n834_adj_814[9]), 
            .I2(n102_c), .I3(n18011), .O(n833_adj_815[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_12 (.CI(n18011), .I0(n834_adj_814[9]), 
            .I1(n102_c), .CO(n18012));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_11_lut (.I0(GND_net), .I1(n834_adj_814[8]), 
            .I2(n102_c), .I3(n18010), .O(n833_adj_815[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_11 (.CI(n18010), .I0(n834_adj_814[8]), 
            .I1(n102_c), .CO(n18011));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_10_lut (.I0(GND_net), .I1(n834_adj_814[7]), 
            .I2(n102_c), .I3(n18009), .O(n833_adj_815[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_10 (.CI(n18009), .I0(n834_adj_814[7]), 
            .I1(n102_c), .CO(n18010));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_9_lut (.I0(GND_net), .I1(n834_adj_814[6]), 
            .I2(n102_c), .I3(n18008), .O(n833_adj_815[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_9 (.CI(n18008), .I0(n834_adj_814[6]), 
            .I1(n102_c), .CO(n18009));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_8_lut (.I0(GND_net), .I1(n834_adj_814[5]), 
            .I2(n102_c), .I3(n18007), .O(n833_adj_815[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_8 (.CI(n18007), .I0(n834_adj_814[5]), 
            .I1(n102_c), .CO(n18008));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_7_lut (.I0(GND_net), .I1(n834_adj_814[4]), 
            .I2(n102_c), .I3(n18006), .O(n833_adj_815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_7 (.CI(n18006), .I0(n834_adj_814[4]), 
            .I1(n102_c), .CO(n18007));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_6_lut (.I0(GND_net), .I1(n834_adj_814[3]), 
            .I2(n102_c), .I3(n18005), .O(n833_adj_815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_6 (.CI(n18005), .I0(n834_adj_814[3]), 
            .I1(n102_c), .CO(n18006));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_5_lut (.I0(GND_net), .I1(n834_adj_814[2]), 
            .I2(n102_c), .I3(n18004), .O(n833_adj_815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_5 (.CI(n18004), .I0(n834_adj_814[2]), 
            .I1(n102_c), .CO(n18005));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_4_lut (.I0(GND_net), .I1(n834_adj_814[1]), 
            .I2(n102_c), .I3(n18003), .O(n833_adj_815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_4 (.CI(n18003), .I0(n834_adj_814[1]), 
            .I1(n102_c), .CO(n18004));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_3_lut (.I0(GND_net), .I1(n834_adj_814[0]), 
            .I2(n102_c), .I3(n18002), .O(n833_adj_815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_3 (.CI(n18002), .I0(n834_adj_814[0]), 
            .I1(n102_c), .CO(n18003));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_2_lut (.I0(GND_net), .I1(n105_c), 
            .I2(n102_c), .I3(GND_net), .O(n833_adj_815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_2 (.CI(GND_net), .I0(n105_c), 
            .I1(n102_c), .CO(n18002));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_16_lut (.I0(GND_net), .I1(n833_adj_815[13]), 
            .I2(n737_c), .I3(n18000), .O(n832_adj_816[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_16 (.CI(n18000), .I0(n833_adj_815[13]), 
            .I1(n737_c), .CO(n739));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_15_lut (.I0(GND_net), .I1(n833_adj_815[12]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17999), .O(Proportional_Gain_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_15 (.CI(n17999), .I0(n833_adj_815[12]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n18000));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_14_lut (.I0(GND_net), .I1(n833_adj_815[11]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17998), .O(Proportional_Gain_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_14 (.CI(n17998), .I0(n833_adj_815[11]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17999));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_13_lut (.I0(GND_net), .I1(n833_adj_815[10]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17997), .O(Proportional_Gain_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_13 (.CI(n17997), .I0(n833_adj_815[10]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17998));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_12_lut (.I0(GND_net), .I1(n833_adj_815[9]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17996), .O(Proportional_Gain_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_12 (.CI(n17996), .I0(n833_adj_815[9]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17997));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_11_lut (.I0(GND_net), .I1(n833_adj_815[8]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17995), .O(Proportional_Gain_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_11 (.CI(n17995), .I0(n833_adj_815[8]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17996));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_10_lut (.I0(GND_net), .I1(n833_adj_815[7]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17994), .O(Proportional_Gain_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_10 (.CI(n17994), .I0(n833_adj_815[7]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17995));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_9_lut (.I0(GND_net), .I1(n833_adj_815[6]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17993), .O(Proportional_Gain_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_9 (.CI(n17993), .I0(n833_adj_815[6]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17994));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_8_lut (.I0(GND_net), .I1(n833_adj_815[5]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17992), .O(Proportional_Gain_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_8 (.CI(n17992), .I0(n833_adj_815[5]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17993));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_7_lut (.I0(GND_net), .I1(n833_adj_815[4]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17991), .O(Proportional_Gain_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_7 (.CI(n17991), .I0(n833_adj_815[4]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17992));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_6_lut (.I0(GND_net), .I1(n833_adj_815[3]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17990), .O(Proportional_Gain_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_6 (.CI(n17990), .I0(n833_adj_815[3]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17991));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_5_lut (.I0(GND_net), .I1(n833_adj_815[2]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17989), .O(Proportional_Gain_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_5 (.CI(n17989), .I0(n833_adj_815[2]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17990));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_4_lut (.I0(GND_net), .I1(n833_adj_815[1]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17988), .O(Proportional_Gain_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_4 (.CI(n17988), .I0(n833_adj_815[1]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17989));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_3_lut (.I0(GND_net), .I1(n833_adj_815[0]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17987), .O(Proportional_Gain_mul_temp[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_3 (.CI(n17987), .I0(n833_adj_815[0]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17988));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_2_lut (.I0(GND_net), .I1(n102_c), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(GND_net), .O(Proportional_Gain_mul_temp[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_2 (.CI(GND_net), .I0(n102_c), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17987));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_8_lut (.I0(GND_net), .I1(n845_adj_818[3]), 
            .I2(n785_c), .I3(n17978), .O(n844_adj_817[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_8 (.CI(n17978), .I0(n845_adj_818[3]), 
            .I1(n785_c), .CO(n787_adj_721));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_7_lut (.I0(GND_net), .I1(n845_adj_818[3]), 
            .I2(n135_c), .I3(n17977), .O(n844_adj_817[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_7 (.CI(n17977), .I0(n845_adj_818[3]), 
            .I1(n135_c), .CO(n17978));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_6_lut (.I0(GND_net), .I1(n845_adj_818[3]), 
            .I2(n135_c), .I3(n17976), .O(n844_adj_817[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_6 (.CI(n17976), .I0(n845_adj_818[3]), 
            .I1(n135_c), .CO(n17977));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_5_lut (.I0(GND_net), .I1(n845_adj_818[2]), 
            .I2(n135_c), .I3(n17975), .O(n844_adj_817[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_5 (.CI(n17975), .I0(n845_adj_818[2]), 
            .I1(n135_c), .CO(n17976));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_4_lut (.I0(GND_net), .I1(n845_adj_818[1]), 
            .I2(n135_c), .I3(n17974), .O(n844_adj_817[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_4 (.CI(n17974), .I0(n845_adj_818[1]), 
            .I1(n135_c), .CO(n17975));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_3_lut (.I0(GND_net), .I1(n845_adj_818[0]), 
            .I2(n135_c), .I3(n17973), .O(n844_adj_817[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_3 (.CI(n17973), .I0(n845_adj_818[0]), 
            .I1(n135_c), .CO(n17974));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_2_lut (.I0(GND_net), .I1(n138_c), 
            .I2(n135_c), .I3(GND_net), .O(n844_adj_817[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_2 (.CI(GND_net), .I0(n138_c), 
            .I1(n135_c), .CO(n17973));
    SB_LUT4 add_4258_17_lut (.I0(GND_net), .I1(n796), .I2(GND_net), .I3(n17972), 
            .O(Proportional_Gain_mul_temp[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4258_16_lut (.I0(GND_net), .I1(n794), .I2(n791_adj_732), 
            .I3(n17971), .O(Proportional_Gain_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_16 (.CI(n17971), .I0(n794), .I1(n791_adj_732), .CO(n17972));
    SB_LUT4 add_4258_15_lut (.I0(GND_net), .I1(n845_adj_818[14]), .I2(n787_adj_721), 
            .I3(n17970), .O(Proportional_Gain_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_15 (.CI(n17970), .I0(n845_adj_818[14]), .I1(n787_adj_721), 
            .CO(n17971));
    SB_LUT4 add_4258_14_lut (.I0(GND_net), .I1(n844_adj_817[14]), .I2(n783_adj_734), 
            .I3(n17969), .O(Proportional_Gain_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_14 (.CI(n17969), .I0(n844_adj_817[14]), .I1(n783_adj_734), 
            .CO(n17970));
    SB_LUT4 add_4258_13_lut (.I0(GND_net), .I1(n843_adj_819[14]), .I2(n779_adj_736), 
            .I3(n17968), .O(Proportional_Gain_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_13 (.CI(n17968), .I0(n843_adj_819[14]), .I1(n779_adj_736), 
            .CO(n17969));
    SB_LUT4 add_4258_12_lut (.I0(GND_net), .I1(n842[14]), .I2(n775), .I3(n17967), 
            .O(Proportional_Gain_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_12 (.CI(n17967), .I0(n842[14]), .I1(n775), .CO(n17968));
    SB_LUT4 add_4258_11_lut (.I0(GND_net), .I1(n841[14]), .I2(n771_adj_598), 
            .I3(n17966), .O(Proportional_Gain_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_11 (.CI(n17966), .I0(n841[14]), .I1(n771_adj_598), 
            .CO(n17967));
    SB_LUT4 add_4258_10_lut (.I0(GND_net), .I1(n840_adj_808[14]), .I2(n767_adj_620), 
            .I3(n17965), .O(Proportional_Gain_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_10 (.CI(n17965), .I0(n840_adj_808[14]), .I1(n767_adj_620), 
            .CO(n17966));
    SB_LUT4 add_4258_9_lut (.I0(GND_net), .I1(n839_adj_809[14]), .I2(n763_adj_636), 
            .I3(n17964), .O(Proportional_Gain_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_9 (.CI(n17964), .I0(n839_adj_809[14]), .I1(n763_adj_636), 
            .CO(n17965));
    SB_LUT4 add_4258_8_lut (.I0(GND_net), .I1(n838_adj_810[14]), .I2(n759_adj_652), 
            .I3(n17963), .O(Proportional_Gain_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_8 (.CI(n17963), .I0(n838_adj_810[14]), .I1(n759_adj_652), 
            .CO(n17964));
    SB_LUT4 add_4258_7_lut (.I0(GND_net), .I1(n837_adj_811[14]), .I2(n755_adj_668), 
            .I3(n17962), .O(Proportional_Gain_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_7 (.CI(n17962), .I0(n837_adj_811[14]), .I1(n755_adj_668), 
            .CO(n17963));
    SB_LUT4 add_4258_6_lut (.I0(GND_net), .I1(n836_adj_812[14]), .I2(n751_adj_684), 
            .I3(n17961), .O(Proportional_Gain_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_6 (.CI(n17961), .I0(n836_adj_812[14]), .I1(n751_adj_684), 
            .CO(n17962));
    SB_LUT4 add_4258_5_lut (.I0(GND_net), .I1(n835_adj_813[14]), .I2(n747_adj_700), 
            .I3(n17960), .O(Proportional_Gain_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_5 (.CI(n17960), .I0(n835_adj_813[14]), .I1(n747_adj_700), 
            .CO(n17961));
    SB_LUT4 add_4258_4_lut (.I0(GND_net), .I1(n834_adj_814[14]), .I2(n743_adj_716), 
            .I3(n17959), .O(Proportional_Gain_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_4 (.CI(n17959), .I0(n834_adj_814[14]), .I1(n743_adj_716), 
            .CO(n17960));
    SB_LUT4 add_4258_3_lut (.I0(GND_net), .I1(n833_adj_815[14]), .I2(n739), 
            .I3(n17958), .O(Proportional_Gain_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_3 (.CI(n17958), .I0(n833_adj_815[14]), .I1(n739), 
            .CO(n17959));
    SB_LUT4 add_4258_2_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(\Error_sub_temp[31] ), 
            .I3(n17957), .O(Proportional_Gain_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4258_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4258_2 (.CI(n17957), .I0(\Product_mul_temp[26] ), .I1(\Error_sub_temp[31] ), 
            .CO(n17958));
    SB_CARRY add_4258_1 (.CI(GND_net), .I0(n832_adj_816[14]), .I1(n832_adj_816[14]), 
            .CO(n17957));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_10_lut (.I0(GND_net), .I1(n844_adj_817[5]), 
            .I2(n781_c), .I3(n17734), .O(n843_adj_819[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_10 (.CI(n17734), .I0(n844_adj_817[5]), 
            .I1(n781_c), .CO(n783_adj_734));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_9_lut (.I0(GND_net), .I1(n844_adj_817[5]), 
            .I2(n132_c), .I3(n17733), .O(n843_adj_819[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_9 (.CI(n17733), .I0(n844_adj_817[5]), 
            .I1(n132_c), .CO(n17734));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_8_lut (.I0(GND_net), .I1(n844_adj_817[5]), 
            .I2(n132_c), .I3(n17732), .O(n843_adj_819[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_8 (.CI(n17661), .I0(n842[5]), 
            .I1(n126_c), .CO(n17662));
    SB_CARRY paramCurrentControlP_15__I_0_add_572_8 (.CI(n17732), .I0(n844_adj_817[5]), 
            .I1(n132_c), .CO(n17733));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_7_lut (.I0(GND_net), .I1(n844_adj_817[4]), 
            .I2(n132_c), .I3(n17731), .O(n843_adj_819[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_7_lut (.I0(GND_net), .I1(n842[4]), 
            .I2(n126_c), .I3(n17660), .O(n841[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_7 (.CI(n17660), .I0(n842[4]), 
            .I1(n126_c), .CO(n17661));
    SB_CARRY paramCurrentControlP_15__I_0_add_572_7 (.CI(n17731), .I0(n844_adj_817[4]), 
            .I1(n132_c), .CO(n17732));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_6_lut (.I0(GND_net), .I1(n842[3]), 
            .I2(n126_c), .I3(n17659), .O(n841[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_6_lut (.I0(GND_net), .I1(n844_adj_817[3]), 
            .I2(n132_c), .I3(n17730), .O(n843_adj_819[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_6 (.CI(n17730), .I0(n844_adj_817[3]), 
            .I1(n132_c), .CO(n17731));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_12_lut (.I0(GND_net), .I1(n843_adj_819[7]), 
            .I2(n777_c), .I3(n17865), .O(n842[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_12 (.CI(n17865), .I0(n843_adj_819[7]), 
            .I1(n777_c), .CO(n779_adj_736));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_11_lut (.I0(GND_net), .I1(n843_adj_819[7]), 
            .I2(n129_c), .I3(n17864), .O(n842[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_11 (.CI(n17864), .I0(n843_adj_819[7]), 
            .I1(n129_c), .CO(n17865));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_10_lut (.I0(GND_net), .I1(n843_adj_819[7]), 
            .I2(n129_c), .I3(n17863), .O(n842[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_10 (.CI(n17863), .I0(n843_adj_819[7]), 
            .I1(n129_c), .CO(n17864));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_9_lut (.I0(GND_net), .I1(n843_adj_819[6]), 
            .I2(n129_c), .I3(n17862), .O(n842[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_9 (.CI(n17862), .I0(n843_adj_819[6]), 
            .I1(n129_c), .CO(n17863));
    SB_LUT4 add_560_33_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[31]), 
            .I3(n15943), .O(Saturate_out1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_32_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[30]), 
            .I3(n15942), .O(\Add_add_temp[34] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_32 (.CI(n15942), .I0(Switch_out1[31]), .I1(currentControlITerm[30]), 
            .CO(n15943));
    SB_LUT4 add_560_31_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[29]), 
            .I3(n15941), .O(\Add_add_temp[33] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_31 (.CI(n15941), .I0(Switch_out1[31]), .I1(currentControlITerm[29]), 
            .CO(n15942));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_8_lut (.I0(GND_net), .I1(n843_adj_819[5]), 
            .I2(n129_c), .I3(n17861), .O(n842[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_560_30_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[28]), 
            .I3(n15940), .O(\Add_add_temp[32] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_30 (.CI(n15940), .I0(Switch_out1[31]), .I1(currentControlITerm[28]), 
            .CO(n15941));
    SB_LUT4 add_560_29_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[27]), 
            .I3(n15939), .O(\Add_add_temp[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_8 (.CI(n17861), .I0(n843_adj_819[5]), 
            .I1(n129_c), .CO(n17862));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_7_lut (.I0(GND_net), .I1(n843_adj_819[4]), 
            .I2(n129_c), .I3(n17860), .O(n842[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_7 (.CI(n17860), .I0(n843_adj_819[4]), 
            .I1(n129_c), .CO(n17861));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_6_lut (.I0(GND_net), .I1(n843_adj_819[3]), 
            .I2(n129_c), .I3(n17859), .O(n842[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_29 (.CI(n15939), .I0(Switch_out1[31]), .I1(currentControlITerm[27]), 
            .CO(n15940));
    SB_LUT4 add_560_28_lut (.I0(GND_net), .I1(Switch_out1[30]), .I2(currentControlITerm[26]), 
            .I3(n15938), .O(\Add_add_temp[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_28 (.CI(n15938), .I0(Switch_out1[30]), .I1(currentControlITerm[26]), 
            .CO(n15939));
    SB_LUT4 add_560_27_lut (.I0(GND_net), .I1(Switch_out1[29]), .I2(currentControlITerm[25]), 
            .I3(n15937), .O(\Add_add_temp[29] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_27 (.CI(n15937), .I0(Switch_out1[29]), .I1(currentControlITerm[25]), 
            .CO(n15938));
    SB_LUT4 add_560_26_lut (.I0(GND_net), .I1(Switch_out1[28]), .I2(currentControlITerm[24]), 
            .I3(n15936), .O(\Add_add_temp[28] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_26 (.CI(n15936), .I0(Switch_out1[28]), .I1(currentControlITerm[24]), 
            .CO(n15937));
    SB_LUT4 add_560_25_lut (.I0(GND_net), .I1(Switch_out1[27]), .I2(currentControlITerm[23]), 
            .I3(n15935), .O(\Add_add_temp[27] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_25 (.CI(n15935), .I0(Switch_out1[27]), .I1(currentControlITerm[23]), 
            .CO(n15936));
    SB_LUT4 add_560_24_lut (.I0(GND_net), .I1(Switch_out1[26]), .I2(currentControlITerm[22]), 
            .I3(n15934), .O(\Add_add_temp[26] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_24 (.CI(n15934), .I0(Switch_out1[26]), .I1(currentControlITerm[22]), 
            .CO(n15935));
    SB_LUT4 add_560_23_lut (.I0(GND_net), .I1(Switch_out1[25]), .I2(currentControlITerm[21]), 
            .I3(n15933), .O(\Add_add_temp[25] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_23 (.CI(n15933), .I0(Switch_out1[25]), .I1(currentControlITerm[21]), 
            .CO(n15934));
    SB_LUT4 add_560_22_lut (.I0(GND_net), .I1(Switch_out1[24]), .I2(currentControlITerm[20]), 
            .I3(n15932), .O(\Add_add_temp[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_22 (.CI(n15932), .I0(Switch_out1[24]), .I1(currentControlITerm[20]), 
            .CO(n15933));
    SB_LUT4 add_560_21_lut (.I0(GND_net), .I1(Switch_out1[23]), .I2(currentControlITerm[19]), 
            .I3(n15931), .O(\Add_add_temp[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_21 (.CI(n15931), .I0(Switch_out1[23]), .I1(currentControlITerm[19]), 
            .CO(n15932));
    SB_LUT4 add_560_20_lut (.I0(GND_net), .I1(Switch_out1[22]), .I2(currentControlITerm[18]), 
            .I3(n15930), .O(\Add_add_temp[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_20 (.CI(n15930), .I0(Switch_out1[22]), .I1(currentControlITerm[18]), 
            .CO(n15931));
    SB_LUT4 add_560_19_lut (.I0(GND_net), .I1(Switch_out1[21]), .I2(currentControlITerm[17]), 
            .I3(n15929), .O(\Add_add_temp[21] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_19 (.CI(n15929), .I0(Switch_out1[21]), .I1(currentControlITerm[17]), 
            .CO(n15930));
    SB_LUT4 add_560_18_lut (.I0(GND_net), .I1(Switch_out1[20]), .I2(currentControlITerm[16]), 
            .I3(n15928), .O(\Add_add_temp[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_18 (.CI(n15928), .I0(Switch_out1[20]), .I1(currentControlITerm[16]), 
            .CO(n15929));
    SB_LUT4 add_560_17_lut (.I0(GND_net), .I1(Switch_out1[19]), .I2(currentControlITerm[15]), 
            .I3(n15927), .O(\Add_add_temp[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_17 (.CI(n15927), .I0(Switch_out1[19]), .I1(currentControlITerm[15]), 
            .CO(n15928));
    SB_LUT4 add_560_16_lut (.I0(GND_net), .I1(Switch_out1[18]), .I2(currentControlITerm[14]), 
            .I3(n15926), .O(\Add_add_temp[18] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_16 (.CI(n15926), .I0(Switch_out1[18]), .I1(currentControlITerm[14]), 
            .CO(n15927));
    SB_LUT4 add_560_15_lut (.I0(GND_net), .I1(Switch_out1[17]), .I2(currentControlITerm[13]), 
            .I3(n15925), .O(\Add_add_temp[17] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_15 (.CI(n15925), .I0(Switch_out1[17]), .I1(currentControlITerm[13]), 
            .CO(n15926));
    SB_LUT4 add_560_14_lut (.I0(GND_net), .I1(Switch_out1[16]), .I2(currentControlITerm[12]), 
            .I3(n15924), .O(\Add_add_temp[16] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_14 (.CI(n15924), .I0(Switch_out1[16]), .I1(currentControlITerm[12]), 
            .CO(n15925));
    SB_LUT4 add_560_13_lut (.I0(GND_net), .I1(Switch_out1[15]), .I2(currentControlITerm[11]), 
            .I3(n15923), .O(\Add_add_temp[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_13 (.CI(n15923), .I0(Switch_out1[15]), .I1(currentControlITerm[11]), 
            .CO(n15924));
    SB_LUT4 add_560_12_lut (.I0(GND_net), .I1(Switch_out1[14]), .I2(currentControlITerm[10]), 
            .I3(n15922), .O(\Add_add_temp[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_12 (.CI(n15922), .I0(Switch_out1[14]), .I1(currentControlITerm[10]), 
            .CO(n15923));
    SB_LUT4 add_560_11_lut (.I0(GND_net), .I1(Switch_out1[13]), .I2(currentControlITerm[9]), 
            .I3(n15921), .O(\Add_add_temp[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_11 (.CI(n15921), .I0(Switch_out1[13]), .I1(currentControlITerm[9]), 
            .CO(n15922));
    SB_LUT4 add_560_10_lut (.I0(GND_net), .I1(Switch_out1[12]), .I2(currentControlITerm[8]), 
            .I3(n15920), .O(\Add_add_temp[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_10 (.CI(n15920), .I0(Switch_out1[12]), .I1(currentControlITerm[8]), 
            .CO(n15921));
    SB_LUT4 add_560_9_lut (.I0(GND_net), .I1(Switch_out1[11]), .I2(preSatVoltage[0]), 
            .I3(n15919), .O(\Add_add_temp[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_9 (.CI(n15919), .I0(Switch_out1[11]), .I1(preSatVoltage[0]), 
            .CO(n15920));
    SB_LUT4 add_560_8_lut (.I0(GND_net), .I1(Switch_out1[10]), .I2(currentControlITerm[6]), 
            .I3(n15918), .O(\Add_add_temp[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_8 (.CI(n15918), .I0(Switch_out1[10]), .I1(currentControlITerm[6]), 
            .CO(n15919));
    SB_LUT4 add_560_7_lut (.I0(GND_net), .I1(Switch_out1[9]), .I2(currentControlITerm[5]), 
            .I3(n15917), .O(\Add_add_temp[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_7 (.CI(n15917), .I0(Switch_out1[9]), .I1(currentControlITerm[5]), 
            .CO(n15918));
    SB_LUT4 add_560_6_lut (.I0(GND_net), .I1(Switch_out1[8]), .I2(currentControlITerm[4]), 
            .I3(n15916), .O(\Add_add_temp[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_6 (.CI(n15916), .I0(Switch_out1[8]), .I1(currentControlITerm[4]), 
            .CO(n15917));
    SB_LUT4 add_560_5_lut (.I0(GND_net), .I1(Switch_out1[7]), .I2(currentControlITerm[3]), 
            .I3(n15915), .O(\Add_add_temp[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_5 (.CI(n15915), .I0(Switch_out1[7]), .I1(currentControlITerm[3]), 
            .CO(n15916));
    SB_LUT4 add_560_4_lut (.I0(GND_net), .I1(Switch_out1[6]), .I2(currentControlITerm[2]), 
            .I3(n15914), .O(\Add_add_temp[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_4 (.CI(n15914), .I0(Switch_out1[6]), .I1(currentControlITerm[2]), 
            .CO(n15915));
    SB_LUT4 add_560_3_lut (.I0(GND_net), .I1(Switch_out1[5]), .I2(currentControlITerm[1]), 
            .I3(n15913), .O(\Add_add_temp[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_3 (.CI(n15913), .I0(Switch_out1[5]), .I1(currentControlITerm[1]), 
            .CO(n15914));
    SB_LUT4 add_560_2_lut (.I0(GND_net), .I1(Switch_out1[4]), .I2(currentControlITerm[0]), 
            .I3(GND_net), .O(\Add_add_temp[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_560_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_560_2 (.CI(GND_net), .I0(Switch_out1[4]), .I1(currentControlITerm[0]), 
            .CO(n15913));
    SB_LUT4 add_548_32_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[30]), 
            .I2(currentControlITerm[31]), .I3(n15912), .O(Voltage_1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_548_31_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[29]), 
            .I2(currentControlITerm[31]), .I3(n15911), .O(preSatVoltage[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_31 (.CI(n15911), .I0(Proportional_Gain_mul_temp[29]), 
            .I1(currentControlITerm[31]), .CO(n15912));
    SB_LUT4 add_548_30_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[28]), 
            .I2(currentControlITerm[31]), .I3(n15910), .O(preSatVoltage[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_30 (.CI(n15910), .I0(Proportional_Gain_mul_temp[28]), 
            .I1(currentControlITerm[31]), .CO(n15911));
    SB_LUT4 add_548_29_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[27]), 
            .I2(currentControlITerm[31]), .I3(n15909), .O(preSatVoltage[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_29 (.CI(n15909), .I0(Proportional_Gain_mul_temp[27]), 
            .I1(currentControlITerm[31]), .CO(n15910));
    SB_LUT4 add_548_28_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[26]), 
            .I2(currentControlITerm[31]), .I3(n15908), .O(preSatVoltage[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_28 (.CI(n15908), .I0(Proportional_Gain_mul_temp[26]), 
            .I1(currentControlITerm[31]), .CO(n15909));
    SB_LUT4 add_548_27_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[25]), 
            .I2(currentControlITerm[31]), .I3(n15907), .O(preSatVoltage[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_27 (.CI(n15907), .I0(Proportional_Gain_mul_temp[25]), 
            .I1(currentControlITerm[31]), .CO(n15908));
    SB_LUT4 add_548_26_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[24]), 
            .I2(currentControlITerm[31]), .I3(n15906), .O(preSatVoltage[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_26 (.CI(n15906), .I0(Proportional_Gain_mul_temp[24]), 
            .I1(currentControlITerm[31]), .CO(n15907));
    SB_LUT4 add_548_25_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[23]), 
            .I2(currentControlITerm[31]), .I3(n15905), .O(preSatVoltage[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_25 (.CI(n15905), .I0(Proportional_Gain_mul_temp[23]), 
            .I1(currentControlITerm[31]), .CO(n15906));
    SB_LUT4 add_548_24_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[22]), 
            .I2(currentControlITerm[30]), .I3(n15904), .O(\preSatVoltage[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_24 (.CI(n15904), .I0(Proportional_Gain_mul_temp[22]), 
            .I1(currentControlITerm[30]), .CO(n15905));
    SB_LUT4 add_548_23_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[21]), 
            .I2(currentControlITerm[29]), .I3(n15903), .O(\preSatVoltage[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_23 (.CI(n15903), .I0(Proportional_Gain_mul_temp[21]), 
            .I1(currentControlITerm[29]), .CO(n15904));
    SB_LUT4 add_548_22_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[20]), 
            .I2(currentControlITerm[28]), .I3(n15902), .O(preSatVoltage[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_22 (.CI(n15902), .I0(Proportional_Gain_mul_temp[20]), 
            .I1(currentControlITerm[28]), .CO(n15903));
    SB_LUT4 add_548_21_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[19]), 
            .I2(currentControlITerm[27]), .I3(n15901), .O(preSatVoltage[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_21 (.CI(n15901), .I0(Proportional_Gain_mul_temp[19]), 
            .I1(currentControlITerm[27]), .CO(n15902));
    SB_LUT4 add_548_20_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[18]), 
            .I2(currentControlITerm[26]), .I3(n15900), .O(\preSatVoltage[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_20 (.CI(n15900), .I0(Proportional_Gain_mul_temp[18]), 
            .I1(currentControlITerm[26]), .CO(n15901));
    SB_LUT4 add_548_19_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[17]), 
            .I2(currentControlITerm[25]), .I3(n15899), .O(preSatVoltage[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_19 (.CI(n15899), .I0(Proportional_Gain_mul_temp[17]), 
            .I1(currentControlITerm[25]), .CO(n15900));
    SB_LUT4 add_548_18_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[16]), 
            .I2(currentControlITerm[24]), .I3(n15898), .O(preSatVoltage[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_18 (.CI(n15898), .I0(Proportional_Gain_mul_temp[16]), 
            .I1(currentControlITerm[24]), .CO(n15899));
    SB_LUT4 add_548_17_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[15]), 
            .I2(currentControlITerm[23]), .I3(n15897), .O(preSatVoltage[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_17 (.CI(n15897), .I0(Proportional_Gain_mul_temp[15]), 
            .I1(currentControlITerm[23]), .CO(n15898));
    SB_LUT4 add_548_16_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[14]), 
            .I2(currentControlITerm[22]), .I3(n15896), .O(preSatVoltage[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_16 (.CI(n15896), .I0(Proportional_Gain_mul_temp[14]), 
            .I1(currentControlITerm[22]), .CO(n15897));
    SB_LUT4 add_548_15_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[13]), 
            .I2(currentControlITerm[21]), .I3(n15895), .O(preSatVoltage[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_15 (.CI(n15895), .I0(Proportional_Gain_mul_temp[13]), 
            .I1(currentControlITerm[21]), .CO(n15896));
    SB_LUT4 add_548_14_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[12]), 
            .I2(currentControlITerm[20]), .I3(n15894), .O(\preSatVoltage[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_14 (.CI(n15894), .I0(Proportional_Gain_mul_temp[12]), 
            .I1(currentControlITerm[20]), .CO(n15895));
    SB_LUT4 add_548_13_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[11]), 
            .I2(currentControlITerm[19]), .I3(n15893), .O(\preSatVoltage[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_13 (.CI(n15893), .I0(Proportional_Gain_mul_temp[11]), 
            .I1(currentControlITerm[19]), .CO(n15894));
    SB_LUT4 add_548_12_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[10]), 
            .I2(currentControlITerm[18]), .I3(n15892), .O(preSatVoltage[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_12 (.CI(n15892), .I0(Proportional_Gain_mul_temp[10]), 
            .I1(currentControlITerm[18]), .CO(n15893));
    SB_LUT4 add_548_11_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[9]), 
            .I2(currentControlITerm[17]), .I3(n15891), .O(\preSatVoltage[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_11 (.CI(n15891), .I0(Proportional_Gain_mul_temp[9]), 
            .I1(currentControlITerm[17]), .CO(n15892));
    SB_LUT4 add_548_10_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[8]), 
            .I2(currentControlITerm[16]), .I3(n15890), .O(preSatVoltage[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_10 (.CI(n15890), .I0(Proportional_Gain_mul_temp[8]), 
            .I1(currentControlITerm[16]), .CO(n15891));
    SB_LUT4 add_548_9_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[7]), 
            .I2(currentControlITerm[15]), .I3(n15889), .O(preSatVoltage[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_9 (.CI(n15889), .I0(Proportional_Gain_mul_temp[7]), 
            .I1(currentControlITerm[15]), .CO(n15890));
    SB_LUT4 add_548_8_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[6]), 
            .I2(currentControlITerm[14]), .I3(n15888), .O(preSatVoltage[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_8 (.CI(n15888), .I0(Proportional_Gain_mul_temp[6]), 
            .I1(currentControlITerm[14]), .CO(n15889));
    SB_LUT4 add_548_7_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[5]), 
            .I2(currentControlITerm[13]), .I3(n15887), .O(preSatVoltage[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_7 (.CI(n15887), .I0(Proportional_Gain_mul_temp[5]), 
            .I1(currentControlITerm[13]), .CO(n15888));
    SB_LUT4 add_548_6_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[4]), 
            .I2(currentControlITerm[12]), .I3(n15886), .O(preSatVoltage[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_6 (.CI(n15886), .I0(Proportional_Gain_mul_temp[4]), 
            .I1(currentControlITerm[12]), .CO(n15887));
    SB_LUT4 add_548_5_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[3]), 
            .I2(currentControlITerm[11]), .I3(n15885), .O(preSatVoltage[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_5 (.CI(n15885), .I0(Proportional_Gain_mul_temp[3]), 
            .I1(currentControlITerm[11]), .CO(n15886));
    SB_LUT4 add_548_4_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[2]), 
            .I2(currentControlITerm[10]), .I3(n15884), .O(preSatVoltage[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_4 (.CI(n15884), .I0(Proportional_Gain_mul_temp[2]), 
            .I1(currentControlITerm[10]), .CO(n15885));
    SB_LUT4 add_548_3_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[1]), 
            .I2(currentControlITerm[9]), .I3(n15883), .O(preSatVoltage[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_548_3 (.CI(n15883), .I0(Proportional_Gain_mul_temp[1]), 
            .I1(currentControlITerm[9]), .CO(n15884));
    SB_LUT4 add_548_2_lut (.I0(preSatVoltage[0]), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(currentControlITerm[8]), .I3(GND_net), .O(n20174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_548_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_548_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(currentControlITerm[8]), .CO(n15883));
    SB_CARRY paramCurrentControlP_15__I_0_add_571_6 (.CI(n17859), .I0(n843_adj_819[3]), 
            .I1(n129_c), .CO(n17860));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_5_lut (.I0(GND_net), .I1(n843_adj_819[2]), 
            .I2(n129_c), .I3(n17858), .O(n842[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_5 (.CI(n17858), .I0(n843_adj_819[2]), 
            .I1(n129_c), .CO(n17859));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_4_lut (.I0(GND_net), .I1(n843_adj_819[1]), 
            .I2(n129_c), .I3(n17857), .O(n842[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_4 (.CI(n17857), .I0(n843_adj_819[1]), 
            .I1(n129_c), .CO(n17858));
    SB_CARRY paramCurrentControlP_15__I_0_add_570_6 (.CI(n17659), .I0(n842[3]), 
            .I1(n126_c), .CO(n17660));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_5_lut (.I0(GND_net), .I1(n842[2]), 
            .I2(n126_c), .I3(n17658), .O(n841[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_3_lut (.I0(GND_net), .I1(n843_adj_819[0]), 
            .I2(n129_c), .I3(n17856), .O(n842[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_3 (.CI(n17856), .I0(n843_adj_819[0]), 
            .I1(n129_c), .CO(n17857));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_2_lut (.I0(GND_net), .I1(n132_c), 
            .I2(n129_c), .I3(GND_net), .O(n842[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_5_lut (.I0(GND_net), .I1(n844_adj_817[2]), 
            .I2(n132_c), .I3(n17729), .O(n843_adj_819[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_2 (.CI(GND_net), .I0(n132_c), 
            .I1(n129_c), .CO(n17856));
    SB_CARRY paramCurrentControlP_15__I_0_add_570_5 (.CI(n17658), .I0(n842[2]), 
            .I1(n126_c), .CO(n17659));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_4_lut (.I0(GND_net), .I1(n842[1]), 
            .I2(n126_c), .I3(n17657), .O(n841[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_5 (.CI(n17729), .I0(n844_adj_817[2]), 
            .I1(n132_c), .CO(n17730));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_4_lut (.I0(GND_net), .I1(n844_adj_817[1]), 
            .I2(n132_c), .I3(n17728), .O(n843_adj_819[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_4 (.CI(n17657), .I0(n842[1]), 
            .I1(n126_c), .CO(n17658));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_3_lut (.I0(GND_net), .I1(n842[0]), 
            .I2(n126_c), .I3(n17656), .O(n841[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_3 (.CI(n17656), .I0(n842[0]), 
            .I1(n126_c), .CO(n17657));
    SB_CARRY paramCurrentControlP_15__I_0_add_572_4 (.CI(n17728), .I0(n844_adj_817[1]), 
            .I1(n132_c), .CO(n17729));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_3_lut (.I0(GND_net), .I1(n844_adj_817[0]), 
            .I2(n132_c), .I3(n17727), .O(n843_adj_819[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_3 (.CI(n17727), .I0(n844_adj_817[0]), 
            .I1(n132_c), .CO(n17728));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_2_lut (.I0(GND_net), .I1(n135_c), 
            .I2(n132_c), .I3(GND_net), .O(n843_adj_819[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_2 (.CI(GND_net), .I0(n135_c), 
            .I1(n132_c), .CO(n17727));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_2_lut (.I0(GND_net), .I1(n129_c), 
            .I2(n126_c), .I3(GND_net), .O(n841[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_2 (.CI(GND_net), .I0(n129_c), 
            .I1(n126_c), .CO(n17656));
    SB_LUT4 add_308_30_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[29]), 
            .I3(n15747), .O(\Error_sub_temp[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_308_29_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[28]), 
            .I3(n15746), .O(\Error_sub_temp[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_29 (.CI(n15746), .I0(\Product_mul_temp[26] ), .I1(n1[28]), 
            .CO(n15747));
    SB_LUT4 add_308_28_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[27]), 
            .I3(n15745), .O(Error_sub_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_28 (.CI(n15745), .I0(\Product_mul_temp[26] ), .I1(n1[27]), 
            .CO(n15746));
    SB_LUT4 add_308_27_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[26]), 
            .I3(n15744), .O(Error_sub_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_27 (.CI(n15744), .I0(\Product_mul_temp[26] ), .I1(n1[26]), 
            .CO(n15745));
    SB_LUT4 add_308_26_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[25]), 
            .I3(n15743), .O(Error_sub_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_26 (.CI(n15743), .I0(\Product_mul_temp[26] ), .I1(n1[25]), 
            .CO(n15744));
    SB_LUT4 add_308_25_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[24]), 
            .I3(n15742), .O(Error_sub_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_25 (.CI(n15742), .I0(\Product_mul_temp[26] ), .I1(n1[24]), 
            .CO(n15743));
    SB_LUT4 add_308_24_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[23]), 
            .I3(n15741), .O(Error_sub_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_24 (.CI(n15741), .I0(\Product_mul_temp[26] ), .I1(n1[23]), 
            .CO(n15742));
    SB_LUT4 add_308_23_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[22]), 
            .I3(n15740), .O(Error_sub_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_23 (.CI(n15740), .I0(\Product_mul_temp[26] ), .I1(n1[22]), 
            .CO(n15741));
    SB_LUT4 add_308_22_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[21]), 
            .I3(n15739), .O(Error_sub_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_22 (.CI(n15739), .I0(\Product_mul_temp[26] ), .I1(n1[21]), 
            .CO(n15740));
    SB_LUT4 add_308_21_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[20]), 
            .I3(n15738), .O(Error_sub_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_21 (.CI(n15738), .I0(\Product_mul_temp[26] ), .I1(n1[20]), 
            .CO(n15739));
    SB_LUT4 add_308_20_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[19]), 
            .I3(n15737), .O(Error_sub_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_20 (.CI(n15737), .I0(\Product_mul_temp[26] ), .I1(n1[19]), 
            .CO(n15738));
    SB_LUT4 add_308_19_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[18]), 
            .I3(n15736), .O(Error_sub_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_19 (.CI(n15736), .I0(\Product_mul_temp[26] ), .I1(n1[18]), 
            .CO(n15737));
    SB_LUT4 add_308_18_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[17]), 
            .I3(n15735), .O(Error_sub_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_18 (.CI(n15735), .I0(\Product_mul_temp[26] ), .I1(n1[17]), 
            .CO(n15736));
    SB_LUT4 add_308_17_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[16]), 
            .I3(n15734), .O(Error_sub_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_17 (.CI(n15734), .I0(\Product_mul_temp[26] ), .I1(n1[16]), 
            .CO(n15735));
    SB_LUT4 add_308_16_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[15]), 
            .I3(n15733), .O(Error_sub_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_16 (.CI(n15733), .I0(\Product_mul_temp[26] ), .I1(n1[15]), 
            .CO(n15734));
    SB_LUT4 add_308_15_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(n1[14]), 
            .I3(n15732), .O(Error_sub_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_308_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_308_15 (.CI(n15732), .I0(\Product_mul_temp[26] ), .I1(n1[14]), 
            .CO(n15733));
    SB_CARRY add_308_14 (.CI(n15731), .I0(\Product_mul_temp[26] ), .I1(n1[13]), 
            .CO(n15732));
    SB_CARRY add_308_13 (.CI(n15730), .I0(GND_net), .I1(n1[12]), .CO(n15731));
    SB_CARRY add_308_12 (.CI(n15729), .I0(GND_net), .I1(n1[11]), .CO(n15730));
    SB_CARRY add_308_11 (.CI(n15728), .I0(GND_net), .I1(n1[10]), .CO(n15729));
    SB_CARRY add_308_10 (.CI(n15727), .I0(GND_net), .I1(n1[9]), .CO(n15728));
    SB_CARRY add_308_9 (.CI(n15726), .I0(GND_net), .I1(n1[8]), .CO(n15727));
    SB_CARRY add_308_8 (.CI(n15725), .I0(GND_net), .I1(n1[7]), .CO(n15726));
    SB_CARRY add_308_7 (.CI(n15724), .I0(GND_net), .I1(n1[6]), .CO(n15725));
    SB_CARRY add_308_6 (.CI(n15723), .I0(GND_net), .I1(n1[5]), .CO(n15724));
    SB_CARRY add_308_5 (.CI(n15722), .I0(GND_net), .I1(n1[4]), .CO(n15723));
    SB_CARRY add_308_4 (.CI(n15721), .I0(GND_net), .I1(n1[3]), .CO(n15722));
    SB_CARRY add_308_3 (.CI(n15720), .I0(GND_net), .I1(n1[2]), .CO(n15721));
    SB_CARRY add_308_2 (.CI(GND_net), .I0(n31), .I1(n1[1]), .CO(n15720));
    SB_LUT4 paramCurrentControlP_15__I_0_i53_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[25]), .I2(GND_net), .I3(GND_net), .O(n126_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i525_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[25]), .I2(GND_net), .I3(GND_net), .O(n773_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i525_2_lut.LUT_INIT = 16'h2222;
    SB_DFF currentControlITerm_i0 (.Q(currentControlITerm[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(n19765));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i4 (.Q(currentControlITerm[4]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14355));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i31 (.Q(currentControlITerm[31]), .C(pin3_clk_16mhz_N_keep), 
           .D(Saturate_out1[31]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 sub_81_inv_0_i2_1_lut (.I0(\qCurrent[3] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[1]));
    defparam sub_81_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i3_1_lut (.I0(\qCurrent[4] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[2]));
    defparam sub_81_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i4_1_lut (.I0(\qCurrent[5] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));
    defparam sub_81_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i5_1_lut (.I0(\qCurrent[6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));
    defparam sub_81_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i6_1_lut (.I0(\qCurrent[7] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));
    defparam sub_81_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i7_1_lut (.I0(\qCurrent[8] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));
    defparam sub_81_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i8_1_lut (.I0(\qCurrent[9] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));
    defparam sub_81_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i9_1_lut (.I0(\qCurrent[10] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));
    defparam sub_81_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i10_1_lut (.I0(\qCurrent[11] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[9]));
    defparam sub_81_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i11_1_lut (.I0(\qCurrent[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[10]));
    defparam sub_81_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i12_1_lut (.I0(\qCurrent[13] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[11]));
    defparam sub_81_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i13_1_lut (.I0(\qCurrent[14] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[12]));
    defparam sub_81_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i14_1_lut (.I0(\qCurrent[15] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[13]));
    defparam sub_81_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i15_1_lut (.I0(\qCurrent[16] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[14]));
    defparam sub_81_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i16_1_lut (.I0(\qCurrent[17] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[15]));
    defparam sub_81_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i17_1_lut (.I0(\qCurrent[18] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[16]));
    defparam sub_81_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i18_1_lut (.I0(\qCurrent[19] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[17]));
    defparam sub_81_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i19_1_lut (.I0(\qCurrent[20] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[18]));
    defparam sub_81_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i20_1_lut (.I0(\qCurrent[21] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[19]));
    defparam sub_81_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i21_1_lut (.I0(\qCurrent[22] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[20]));
    defparam sub_81_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i22_1_lut (.I0(\qCurrent[23] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[21]));
    defparam sub_81_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i23_1_lut (.I0(\qCurrent[24] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[22]));
    defparam sub_81_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i24_1_lut (.I0(\qCurrent[25] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[23]));
    defparam sub_81_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i25_1_lut (.I0(\qCurrent[26] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[24]));
    defparam sub_81_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i26_1_lut (.I0(\qCurrent[27] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[25]));
    defparam sub_81_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i27_1_lut (.I0(\qCurrent[28] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[26]));
    defparam sub_81_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i28_1_lut (.I0(\qCurrent[29] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[27]));
    defparam sub_81_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i29_1_lut (.I0(\qCurrent[30] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[28]));
    defparam sub_81_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_81_inv_0_i30_1_lut (.I0(\qCurrent[31] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[29]));
    defparam sub_81_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_271 (.I0(n138_c), .I1(n142), .I2(n10_adj_755), 
            .I3(n14_adj_756), .O(n4_adj_757));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_adj_271.LUT_INIT = 16'heca8;
    SB_LUT4 i1_4_lut_adj_272 (.I0(n138_c), .I1(n142), .I2(n14_adj_756), 
            .I3(n10_adj_755), .O(n18_adj_758));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_adj_272.LUT_INIT = 16'heca8;
    SB_LUT4 i2_4_lut (.I0(n142), .I1(n4_adj_757), .I2(n138_c), .I3(n10_adj_755), 
            .O(n19841));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i1_4_lut_adj_273 (.I0(n138_c), .I1(n142), .I2(n19841), .I3(n18_adj_758), 
            .O(n26_adj_759));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_adj_273.LUT_INIT = 16'heca8;
    SB_LUT4 i1_4_lut_adj_274 (.I0(n138_c), .I1(n7_adj_760), .I2(Error_sub_temp[29]), 
            .I3(n26_adj_759), .O(n791_adj_732));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_adj_274.LUT_INIT = 16'hcecc;
    SB_LUT4 i12078_3_lut (.I0(\Product_mul_temp[26] ), .I1(\Error_sub_temp[30] ), 
            .I2(Error_sub_temp[29]), .I3(GND_net), .O(n845_adj_818[0]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i12078_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i2_4_lut_adj_275 (.I0(n141), .I1(n138_c), .I2(Error_sub_temp[29]), 
            .I3(n146), .O(n845_adj_818[1]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_4_lut_adj_275.LUT_INIT = 16'h39c6;
    SB_LUT4 i12085_4_lut (.I0(Error_sub_temp[29]), .I1(n138_c), .I2(n141), 
            .I3(\Error_sub_temp[30] ), .O(n4_adj_761));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i12085_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 i1_2_lut (.I0(\Add_add_temp[5] ), .I1(\Add_add_temp[4] ), .I2(GND_net), 
            .I3(GND_net), .O(n20722));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_276 (.I0(\Add_add_temp[7] ), .I1(\Add_add_temp[8] ), 
            .I2(\Add_add_temp[6] ), .I3(n20722), .O(n19761));
    defparam i1_4_lut_adj_276.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_277 (.I0(\Add_add_temp[11] ), .I1(n19761), .I2(\Add_add_temp[10] ), 
            .I3(\Add_add_temp[9] ), .O(n20704));
    defparam i1_4_lut_adj_277.LUT_INIT = 16'hfaea;
    SB_LUT4 i13263_4_lut (.I0(\Add_add_temp[12] ), .I1(\Add_add_temp[14] ), 
            .I2(\Add_add_temp[13] ), .I3(n20704), .O(n15200));
    defparam i13263_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i6661_2_lut (.I0(n833[13]), .I1(\Error_sub_temp[31] ), .I2(GND_net), 
            .I3(GND_net), .O(n832[14]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(92[30:64])
    defparam i6661_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6663_2_lut (.I0(n833[13]), .I1(\Error_sub_temp[31] ), .I2(GND_net), 
            .I3(GND_net), .O(n8356));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(92[30:64])
    defparam i6663_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_278 (.I0(\Add_add_temp[17] ), .I1(n15200), .I2(\Add_add_temp[16] ), 
            .I3(\Add_add_temp[15] ), .O(n20680));
    defparam i1_4_lut_adj_278.LUT_INIT = 16'hfaea;
    SB_LUT4 i1_4_lut_adj_279 (.I0(\Add_add_temp[19] ), .I1(\Add_add_temp[20] ), 
            .I2(\Add_add_temp[18] ), .I3(n20680), .O(n19733));
    defparam i1_4_lut_adj_279.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_280 (.I0(\Add_add_temp[23] ), .I1(n19733), .I2(\Add_add_temp[22] ), 
            .I3(\Add_add_temp[21] ), .O(n20660));
    defparam i1_4_lut_adj_280.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_281 (.I0(\Add_add_temp[26] ), .I1(n20660), .I2(\Add_add_temp[25] ), 
            .I3(\Add_add_temp[24] ), .O(n20654));
    defparam i1_4_lut_adj_281.LUT_INIT = 16'hfaea;
    SB_LUT4 i1_4_lut_adj_282 (.I0(\Add_add_temp[29] ), .I1(n20654), .I2(\Add_add_temp[28] ), 
            .I3(\Add_add_temp[27] ), .O(n20640));
    defparam i1_4_lut_adj_282.LUT_INIT = 16'hfaea;
    SB_LUT4 i14382_4_lut (.I0(\Add_add_temp[30] ), .I1(\Add_add_temp[32] ), 
            .I2(\Add_add_temp[31] ), .I3(n20640), .O(n19308));
    defparam i14382_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut_adj_283 (.I0(\Add_add_temp[34] ), .I1(Saturate_out1[31]), 
            .I2(\Add_add_temp[33] ), .I3(n19308), .O(Saturate_out1_31__N_267));
    defparam i1_4_lut_adj_283.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_284 (.I0(\Add_add_temp[7] ), .I1(\Add_add_temp[8] ), 
            .I2(\Add_add_temp[6] ), .I3(\Add_add_temp[5] ), .O(n19755));
    defparam i1_4_lut_adj_284.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_285 (.I0(\Add_add_temp[11] ), .I1(n19755), .I2(\Add_add_temp[10] ), 
            .I3(\Add_add_temp[9] ), .O(n20718));
    defparam i1_4_lut_adj_285.LUT_INIT = 16'ha8a0;
    SB_LUT4 i772_4_lut (.I0(\Add_add_temp[12] ), .I1(\Add_add_temp[14] ), 
            .I2(\Add_add_temp[13] ), .I3(n20718), .O(n22_adj_762));
    defparam i772_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_286 (.I0(\Add_add_temp[17] ), .I1(n22_adj_762), 
            .I2(\Add_add_temp[16] ), .I3(\Add_add_temp[15] ), .O(n20694));
    defparam i1_4_lut_adj_286.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_287 (.I0(\Add_add_temp[19] ), .I1(\Add_add_temp[20] ), 
            .I2(\Add_add_temp[18] ), .I3(n20694), .O(n19729));
    defparam i1_4_lut_adj_287.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_3_lut_4_lut (.I0(n142), .I1(\Product_mul_temp[26] ), 
            .I2(Error_sub_temp[29]), .I3(n4_adj_761), .O(n10_adj_755));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_4_lut_4_lut (.I0(\Product_mul_temp[26] ), .I1(Error_sub_temp[29]), 
            .I2(n142), .I3(n26_adj_759), .O(n845_adj_818[14]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h2a52;
    SB_LUT4 i1_4_lut_adj_288 (.I0(\Add_add_temp[23] ), .I1(n19729), .I2(\Add_add_temp[22] ), 
            .I3(\Add_add_temp[21] ), .O(n20676));
    defparam i1_4_lut_adj_288.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Product_mul_temp[26] ), .I1(Error_sub_temp[29]), 
            .I2(n142), .I3(n4_adj_761), .O(n845_adj_818[3]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h80f8;
    SB_LUT4 i2_3_lut_4_lut (.I0(n4_adj_761), .I1(\Product_mul_temp[26] ), 
            .I2(Error_sub_temp[29]), .I3(n142), .O(n845_adj_818[2]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 i1_4_lut_adj_289 (.I0(\Add_add_temp[26] ), .I1(n20676), .I2(\Add_add_temp[25] ), 
            .I3(\Add_add_temp[24] ), .O(n20664));
    defparam i1_4_lut_adj_289.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_290 (.I0(\Add_add_temp[29] ), .I1(n20664), .I2(\Add_add_temp[28] ), 
            .I3(\Add_add_temp[27] ), .O(n20650));
    defparam i1_4_lut_adj_290.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_3_lut_4_lut_adj_291 (.I0(n146), .I1(n141), .I2(n26_adj_759), 
            .I3(\Product_mul_temp[26] ), .O(n7_adj_760));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_3_lut_4_lut_adj_291.LUT_INIT = 16'heee0;
    SB_LUT4 i790_4_lut (.I0(\Add_add_temp[30] ), .I1(\Add_add_temp[32] ), 
            .I2(\Add_add_temp[31] ), .I3(n20650), .O(n58));
    defparam i790_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_4_lut_adj_292 (.I0(\Product_mul_temp[26] ), .I1(Error_sub_temp[29]), 
            .I2(n6_adj_763), .I3(n10_adj_755), .O(n14_adj_756));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_3_lut_4_lut_adj_292.LUT_INIT = 16'hf8f0;
    SB_LUT4 i1_4_lut_adj_293 (.I0(\Add_add_temp[34] ), .I1(Saturate_out1[31]), 
            .I2(\Add_add_temp[33] ), .I3(n58), .O(Saturate_out1_31__N_266));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(121[27:75])
    defparam i1_4_lut_adj_293.LUT_INIT = 16'h2000;
    SB_LUT4 sub_81_inv_0_i1_1_lut_2_lut (.I0(\Product_mul_temp[26] ), .I1(Look_Up_Table_out1_1[0]), 
            .I2(GND_net), .I3(GND_net), .O(n31));
    defparam sub_81_inv_0_i1_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_3_lut_3_lut_4_lut (.I0(n142), .I1(\Product_mul_temp[26] ), 
            .I2(Error_sub_temp[29]), .I3(n4_adj_761), .O(n6_adj_763));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_3_lut_3_lut_4_lut.LUT_INIT = 16'haa80;
    Saturate_Output u_Saturate_Output (.\preSatVoltage[20] (preSatVoltage[20]), 
            .Out_31__N_333(Out_31__N_333), .Out_31__N_332(Out_31__N_332), 
            .Look_Up_Table_out1_1({Look_Up_Table_out1_1}), .n579(n579), 
            .\preSatVoltage[9] (preSatVoltage[9]), .n17(n17), .\preSatVoltage[14] (preSatVoltage[14]), 
            .n267(n267), .\preSatVoltage[11] (preSatVoltage[11]), .n120(n120), 
            .n14(n14), .\preSatVoltage[17] (preSatVoltage[17]), .n414(n414), 
            .n11(n11), .\preSatVoltage[24] (preSatVoltage[24]), .n19604(n19604), 
            .n789(n789), .n785(n785), .n781(n781), .n8(n8), .n777(n777), 
            .n19351(n19351), .n773(n773), .n769(n769), .n765(n765), 
            .n270(n270), .n123(n123), .n761(n761), .n757(n757), .n417(n417), 
            .n753(n753), .n749(n749), .n745(n745), .n741(n741), .n737(n737), 
            .\preSatVoltage[18] (preSatVoltage[18]), .\Product_mul_temp[26] (\Product_mul_temp[26] ), 
            .n489(n489), .\qVoltage[9] (\qVoltage[9] ), .GND_net(GND_net), 
            .n489_adj_19(n489_adj_25), .\preSatVoltage[15] (preSatVoltage[15]), 
            .n342(n342), .\qVoltage[6] (\qVoltage[6] ), .n342_adj_20(n342_adj_26), 
            .\qVoltage[5] (\qVoltage[5] ), .n246(n246), .n288(n288), .n285(n285), 
            .n282(n282), .n279(n279), .n276(n276), .n273(n273), .\qVoltage[15] (\qVoltage[15] ), 
            .n258(n258), .n255(n255), .n252(n252), .n261(n261), .n249(n249), 
            .n44(n44), .n126(n126), .n420(n420), .n129(n129), .n423(n423), 
            .n41(n41), .\preSatVoltage[10] (\preSatVoltage[10] ), .n86(n86), 
            .n89(n89), .n86_adj_21(n86_adj_27), .n83(n83), .n80(n80), 
            .n19702(n19702), .n77(n77), .n74(n74), .n38(n38), .n71(n71), 
            .n68(n68), .n65(n65), .n62(n62), .n59(n59), .n56(n56), 
            .n50(n50), .n53(n53), .n92(n92), .\preSatVoltage[13] (\preSatVoltage[13] ), 
            .n244(n244), .n35(n35), .\qVoltage[4] (\qVoltage[4] ), .\preSatVoltage[12] (\preSatVoltage[12] ), 
            .n195(n195), .\qVoltage[3] (\qVoltage[3] ), .n114(n114), .\qVoltage[2] (\qVoltage[2] ), 
            .n108(n108), .n102(n102), .n99(n99), .\Product2_mul_temp[2] (\Product2_mul_temp[2] ), 
            .n141(n141_adj_28), .n105(n105), .n138(n138), .n135(n135), 
            .n132(n132), .n111(n111), .n32(n32), .\preSatVoltage[19] (\preSatVoltage[19] ), 
            .\qVoltage[10] (\qVoltage[10] ), .n538(n538), .n29(n29), .\preSatVoltage[16] (preSatVoltage[16]), 
            .\preSatVoltage[22] (\preSatVoltage[22] ), .\preSatVoltage[21] (preSatVoltage[21]), 
            .\preSatVoltage[25] (preSatVoltage[25]), .\preSatVoltage[23] (\preSatVoltage[23] ), 
            .\preSatVoltage[28] (preSatVoltage[28]), .\preSatVoltage[27] (preSatVoltage[27]), 
            .\preSatVoltage[26] (preSatVoltage[26]), .\preSatVoltage[29] (preSatVoltage[29]), 
            .\Voltage_1[31] (Voltage_1[31]), .\preSatVoltage[30] (preSatVoltage[30]), 
            .\preSatVoltage[5] (preSatVoltage[5]), .\preSatVoltage[6] (preSatVoltage[6]), 
            .\preSatVoltage[4] (preSatVoltage[4]), .\preSatVoltage[2] (preSatVoltage[2]), 
            .\preSatVoltage[7] (preSatVoltage[7]), .\preSatVoltage[3] (preSatVoltage[3]), 
            .n20174(n20174), .\preSatVoltage[8] (preSatVoltage[8]), .n426(n426), 
            .\qVoltage[13] (\qVoltage[13] ), .n685(n685), .n402(n402), 
            .n429(n429), .n432(n432), .n26(n26), .n391(n391), .n23(n23), 
            .\qVoltage[7] (\qVoltage[7] ), .n391_adj_22(n391_adj_29), .n21(n21), 
            .n576(n576), .n576_adj_23(n576_adj_30), .n573(n573), .n570(n570), 
            .n567(n567), .\qVoltage[12] (\qVoltage[12] ), .n564(n564), 
            .n405(n405), .n628(n628), .n625(n625), .n622(n622), .n435(n435), 
            .n619(n619), .n616(n616), .n613(n613), .n610(n610), .n607(n607), 
            .n601(n601), .n561(n561), .n598(n598), .n595(n595), .n592(n592), 
            .n589(n589), .n604(n604), .n631(n631), .\qVoltage[8] (\qVoltage[8] ), 
            .n558(n558), .n20(n20), .n264(n264), .n117(n117), .n411(n411), 
            .n587(n587), .n587_adj_24(n587_adj_31), .n582(n582), .n393(n393), 
            .n408(n408), .n555(n555), .n552(n552), .n549(n549), .n396(n396), 
            .n399(n399), .n546(n546), .\qVoltage[14] (\qVoltage[14] ), 
            .n543(n543), .n540(n540)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(148[19] 150[39])
    
endmodule
//
// Verilog Description of module Saturate_Output
//

module Saturate_Output (\preSatVoltage[20] , Out_31__N_333, Out_31__N_332, 
            Look_Up_Table_out1_1, n579, \preSatVoltage[9] , n17, \preSatVoltage[14] , 
            n267, \preSatVoltage[11] , n120, n14, \preSatVoltage[17] , 
            n414, n11, \preSatVoltage[24] , n19604, n789, n785, 
            n781, n8, n777, n19351, n773, n769, n765, n270, 
            n123, n761, n757, n417, n753, n749, n745, n741, 
            n737, \preSatVoltage[18] , \Product_mul_temp[26] , n489, 
            \qVoltage[9] , GND_net, n489_adj_19, \preSatVoltage[15] , 
            n342, \qVoltage[6] , n342_adj_20, \qVoltage[5] , n246, 
            n288, n285, n282, n279, n276, n273, \qVoltage[15] , 
            n258, n255, n252, n261, n249, n44, n126, n420, n129, 
            n423, n41, \preSatVoltage[10] , n86, n89, n86_adj_21, 
            n83, n80, n19702, n77, n74, n38, n71, n68, n65, 
            n62, n59, n56, n50, n53, n92, \preSatVoltage[13] , 
            n244, n35, \qVoltage[4] , \preSatVoltage[12] , n195, \qVoltage[3] , 
            n114, \qVoltage[2] , n108, n102, n99, \Product2_mul_temp[2] , 
            n141, n105, n138, n135, n132, n111, n32, \preSatVoltage[19] , 
            \qVoltage[10] , n538, n29, \preSatVoltage[16] , \preSatVoltage[22] , 
            \preSatVoltage[21] , \preSatVoltage[25] , \preSatVoltage[23] , 
            \preSatVoltage[28] , \preSatVoltage[27] , \preSatVoltage[26] , 
            \preSatVoltage[29] , \Voltage_1[31] , \preSatVoltage[30] , 
            \preSatVoltage[5] , \preSatVoltage[6] , \preSatVoltage[4] , 
            \preSatVoltage[2] , \preSatVoltage[7] , \preSatVoltage[3] , 
            n20174, \preSatVoltage[8] , n426, \qVoltage[13] , n685, 
            n402, n429, n432, n26, n391, n23, \qVoltage[7] , n391_adj_22, 
            n21, n576, n576_adj_23, n573, n570, n567, \qVoltage[12] , 
            n564, n405, n628, n625, n622, n435, n619, n616, 
            n613, n610, n607, n601, n561, n598, n595, n592, 
            n589, n604, n631, \qVoltage[8] , n558, n20, n264, 
            n117, n411, n587, n587_adj_24, n582, n393, n408, n555, 
            n552, n549, n396, n399, n546, \qVoltage[14] , n543, 
            n540) /* synthesis syn_module_defined=1 */ ;
    input \preSatVoltage[20] ;
    output Out_31__N_333;
    output Out_31__N_332;
    input [15:0]Look_Up_Table_out1_1;
    output n579;
    input \preSatVoltage[9] ;
    output n17;
    input \preSatVoltage[14] ;
    output n267;
    input \preSatVoltage[11] ;
    output n120;
    output n14;
    input \preSatVoltage[17] ;
    output n414;
    output n11;
    input \preSatVoltage[24] ;
    output n19604;
    output n789;
    output n785;
    output n781;
    output n8;
    output n777;
    output n19351;
    output n773;
    output n769;
    output n765;
    output n270;
    output n123;
    output n761;
    output n757;
    output n417;
    output n753;
    output n749;
    output n745;
    output n741;
    output n737;
    input \preSatVoltage[18] ;
    input \Product_mul_temp[26] ;
    output n489;
    output \qVoltage[9] ;
    input GND_net;
    output n489_adj_19;
    input \preSatVoltage[15] ;
    output n342;
    output \qVoltage[6] ;
    output n342_adj_20;
    output \qVoltage[5] ;
    output n246;
    output n288;
    output n285;
    output n282;
    output n279;
    output n276;
    output n273;
    output \qVoltage[15] ;
    output n258;
    output n255;
    output n252;
    output n261;
    output n249;
    output n44;
    output n126;
    output n420;
    output n129;
    output n423;
    output n41;
    input \preSatVoltage[10] ;
    output n86;
    output n89;
    output n86_adj_21;
    output n83;
    output n80;
    output n19702;
    output n77;
    output n74;
    output n38;
    output n71;
    output n68;
    output n65;
    output n62;
    output n59;
    output n56;
    output n50;
    output n53;
    output n92;
    input \preSatVoltage[13] ;
    output n244;
    output n35;
    output \qVoltage[4] ;
    input \preSatVoltage[12] ;
    output n195;
    output \qVoltage[3] ;
    output n114;
    output \qVoltage[2] ;
    output n108;
    output n102;
    output n99;
    output \Product2_mul_temp[2] ;
    output n141;
    output n105;
    output n138;
    output n135;
    output n132;
    output n111;
    output n32;
    input \preSatVoltage[19] ;
    output \qVoltage[10] ;
    output n538;
    output n29;
    input \preSatVoltage[16] ;
    input \preSatVoltage[22] ;
    input \preSatVoltage[21] ;
    input \preSatVoltage[25] ;
    input \preSatVoltage[23] ;
    input \preSatVoltage[28] ;
    input \preSatVoltage[27] ;
    input \preSatVoltage[26] ;
    input \preSatVoltage[29] ;
    input \Voltage_1[31] ;
    input \preSatVoltage[30] ;
    input \preSatVoltage[5] ;
    input \preSatVoltage[6] ;
    input \preSatVoltage[4] ;
    input \preSatVoltage[2] ;
    input \preSatVoltage[7] ;
    input \preSatVoltage[3] ;
    input n20174;
    input \preSatVoltage[8] ;
    output n426;
    output \qVoltage[13] ;
    output n685;
    output n402;
    output n429;
    output n432;
    output n26;
    output n391;
    output n23;
    output \qVoltage[7] ;
    output n391_adj_22;
    output n21;
    output n576;
    output n576_adj_23;
    output n573;
    output n570;
    output n567;
    output \qVoltage[12] ;
    output n564;
    output n405;
    output n628;
    output n625;
    output n622;
    output n435;
    output n619;
    output n616;
    output n613;
    output n610;
    output n607;
    output n601;
    output n561;
    output n598;
    output n595;
    output n592;
    output n589;
    output n604;
    output n631;
    output \qVoltage[8] ;
    output n558;
    output n20;
    output n264;
    output n117;
    output n411;
    output n587;
    output n587_adj_24;
    output n582;
    output n393;
    output n408;
    output n555;
    output n552;
    output n549;
    output n396;
    output n399;
    output n546;
    output \qVoltage[14] ;
    output n543;
    output n540;
    
    
    wire n19812, n19827, n20102, n20086, n19890, n19896, n19741, 
        n20180, n22, n19450, n19743, n20108, n20092, n19914, n19920;
    
    SB_LUT4 Q_15__I_0_i391_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[13]), .O(n579));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i391_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i3_4_lut (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), .I2(Out_31__N_333), 
            .I3(Look_Up_Table_out1_1[5]), .O(n17));
    defparam i3_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[7]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[14] ), .O(n267));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_148 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[7]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n120));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_148.LUT_INIT = 16'h4440;
    SB_LUT4 i3_4_lut_adj_149 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[4]), .O(n14));
    defparam i3_4_lut_adj_149.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_150 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[7]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n414));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_150.LUT_INIT = 16'h4440;
    SB_LUT4 i3_4_lut_adj_151 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[3]), .O(n11));
    defparam i3_4_lut_adj_151.LUT_INIT = 16'h0400;
    SB_LUT4 i1_3_lut_4_lut (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), .O(n19604));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_152 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n789));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_152.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_153 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), .O(n785));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_153.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_154 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n781));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_154.LUT_INIT = 16'h000e;
    SB_LUT4 i3_4_lut_adj_155 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[2]), .O(n8));
    defparam i3_4_lut_adj_155.LUT_INIT = 16'h0400;
    SB_LUT4 i1_3_lut_4_lut_adj_156 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), .O(n777));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_156.LUT_INIT = 16'h000e;
    SB_LUT4 i1_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), .I2(\preSatVoltage[9] ), 
            .I3(Look_Up_Table_out1_1[1]), .O(n19351));
    defparam i1_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_3_lut_4_lut_adj_157 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), .O(n773));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_157.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_158 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[8]), .I3(Out_31__N_332), .O(n769));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_158.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_159 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), .O(n765));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_159.LUT_INIT = 16'h000e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_160 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[8]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[14] ), .O(n270));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_160.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_161 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[8]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n123));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_161.LUT_INIT = 16'h4440;
    SB_LUT4 i1_3_lut_4_lut_adj_162 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[6]), .I3(Out_31__N_332), .O(n761));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_162.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_163 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n757));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_163.LUT_INIT = 16'h000e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_164 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[8]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n417));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_164.LUT_INIT = 16'h4440;
    SB_LUT4 i1_3_lut_4_lut_adj_165 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n753));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_165.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_166 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n749));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_166.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_167 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n745));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_167.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_168 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n741));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_168.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_169 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n737));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_169.LUT_INIT = 16'h000e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_170 (.I0(\preSatVoltage[18] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n489));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_170.LUT_INIT = 16'h00d0;
    SB_LUT4 i13211_2_lut_3_lut (.I0(\preSatVoltage[18] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[9] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13211_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_171 (.I0(\preSatVoltage[18] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n489_adj_19));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_171.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_172 (.I0(\preSatVoltage[15] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n342));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_172.LUT_INIT = 16'h00d0;
    SB_LUT4 i13208_2_lut_3_lut (.I0(\preSatVoltage[15] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[6] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13208_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_173 (.I0(\preSatVoltage[15] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n342_adj_20));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_173.LUT_INIT = 16'h00d0;
    SB_LUT4 i13207_2_lut_3_lut (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[5] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13207_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_174 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n246));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_174.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_175 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), .O(n288));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_175.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_176 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n285));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_176.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_177 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), .O(n282));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_177.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_178 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n279));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_178.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_179 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), .O(n276));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_179.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_180 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), .O(n273));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_180.LUT_INIT = 16'h00e0;
    SB_LUT4 i13217_2_lut_3_lut (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[15] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13217_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_181 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n258));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_181.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_182 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n255));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_182.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_183 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n252));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_183.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_184 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n261));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_184.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_185 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n249));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_185.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_186 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[14]), .O(n44));
    defparam i3_4_lut_adj_186.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_187 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[9]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n126));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_187.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_188 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[9]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n420));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_188.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_189 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[10]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n129));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_189.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_190 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[10]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n423));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_190.LUT_INIT = 16'h4440;
    SB_LUT4 i3_4_lut_adj_191 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[13]), .O(n41));
    defparam i3_4_lut_adj_191.LUT_INIT = 16'h0400;
    SB_LUT4 Q_15__I_0_11_i39_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(\Product_mul_temp[26] ), .O(n86));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_11_i39_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i61_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[13]), .O(n89));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i61_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i59_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[12]), .O(n86_adj_21));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i59_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i57_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[11]), .O(n83));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i57_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i55_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[10]), .O(n80));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i55_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_3_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), .I2(\preSatVoltage[9] ), 
            .I3(GND_net), .O(n19702));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 Q_15__I_0_i53_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[9]), .O(n77));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i53_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i51_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[8]), .O(n74));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i51_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_adj_192 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[12]), .O(n38));
    defparam i3_4_lut_adj_192.LUT_INIT = 16'h0400;
    SB_LUT4 Q_15__I_0_i49_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[7]), .O(n71));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i49_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i47_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[6]), .O(n68));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i47_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i45_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[5]), .O(n65));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i45_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i43_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[4]), .O(n62));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i43_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i41_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[3]), .O(n59));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i41_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i39_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[2]), .O(n56));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i39_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i35_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[0]), .O(n50));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i35_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i37_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[1]), .O(n53));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i37_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 Q_15__I_0_i63_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[14]), .O(n92));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam Q_15__I_0_i63_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_193 (.I0(\preSatVoltage[13] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n244));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_193.LUT_INIT = 16'h00d0;
    SB_LUT4 i3_4_lut_adj_194 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[11]), .O(n35));
    defparam i3_4_lut_adj_194.LUT_INIT = 16'h0400;
    SB_LUT4 i13206_2_lut_3_lut (.I0(\preSatVoltage[13] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[4] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13206_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_195 (.I0(\preSatVoltage[12] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n195));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_195.LUT_INIT = 16'h00d0;
    SB_LUT4 i13205_2_lut_3_lut (.I0(\preSatVoltage[12] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[3] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13205_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_196 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n114));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_196.LUT_INIT = 16'h00e0;
    SB_LUT4 i13204_2_lut_3_lut (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[2] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13204_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_197 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n108));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_197.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_198 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n102));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_198.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_199 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n99));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_199.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_200 (.I0(Out_31__N_332), .I1(Out_31__N_333), .I2(\preSatVoltage[9] ), 
            .I3(\Product_mul_temp[26] ), .O(\Product2_mul_temp[2] ));
    defparam i3_4_lut_adj_200.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_201 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), .O(n141));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_201.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_202 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n105));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_202.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_203 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n138));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_203.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_204 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), .O(n135));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_204.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_205 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n132));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_205.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_206 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n111));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_206.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_207 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[10]), .O(n32));
    defparam i3_4_lut_adj_207.LUT_INIT = 16'h0400;
    SB_LUT4 i13212_2_lut_3_lut (.I0(\preSatVoltage[19] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[10] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13212_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_208 (.I0(\preSatVoltage[19] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n538));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_208.LUT_INIT = 16'h00d0;
    SB_LUT4 i3_4_lut_adj_209 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[9]), .O(n29));
    defparam i3_4_lut_adj_209.LUT_INIT = 16'h0400;
    SB_LUT4 i1_4_lut_adj_210 (.I0(\preSatVoltage[12] ), .I1(\preSatVoltage[13] ), 
            .I2(\preSatVoltage[10] ), .I3(\preSatVoltage[11] ), .O(n19812));
    defparam i1_4_lut_adj_210.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_211 (.I0(\preSatVoltage[15] ), .I1(\preSatVoltage[16] ), 
            .I2(n19812), .I3(\preSatVoltage[14] ), .O(n19827));
    defparam i1_4_lut_adj_211.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_212 (.I0(\preSatVoltage[19] ), .I1(\preSatVoltage[18] ), 
            .I2(n19827), .I3(\preSatVoltage[17] ), .O(n20102));
    defparam i1_4_lut_adj_212.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_213 (.I0(\preSatVoltage[22] ), .I1(n20102), .I2(\preSatVoltage[21] ), 
            .I3(\preSatVoltage[20] ), .O(n20086));
    defparam i1_4_lut_adj_213.LUT_INIT = 16'hfaea;
    SB_LUT4 i1_4_lut_adj_214 (.I0(\preSatVoltage[25] ), .I1(\preSatVoltage[24] ), 
            .I2(n20086), .I3(\preSatVoltage[23] ), .O(n19890));
    defparam i1_4_lut_adj_214.LUT_INIT = 16'h8880;
    SB_LUT4 i1_4_lut_adj_215 (.I0(\preSatVoltage[28] ), .I1(\preSatVoltage[27] ), 
            .I2(\preSatVoltage[26] ), .I3(n19890), .O(n19896));
    defparam i1_4_lut_adj_215.LUT_INIT = 16'h8000;
    SB_LUT4 i1223_rep_3_4_lut (.I0(\preSatVoltage[29] ), .I1(\Voltage_1[31] ), 
            .I2(\preSatVoltage[30] ), .I3(n19896), .O(Out_31__N_333));
    defparam i1223_rep_3_4_lut.LUT_INIT = 16'h4ccc;
    SB_LUT4 i1_4_lut_adj_216 (.I0(\preSatVoltage[5] ), .I1(\preSatVoltage[6] ), 
            .I2(\preSatVoltage[4] ), .I3(\preSatVoltage[2] ), .O(n19741));
    defparam i1_4_lut_adj_216.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_217 (.I0(n19741), .I1(\preSatVoltage[7] ), .I2(\preSatVoltage[3] ), 
            .I3(n20174), .O(n20180));
    defparam i1_4_lut_adj_217.LUT_INIT = 16'hfffe;
    SB_LUT4 i1213_4_lut (.I0(\preSatVoltage[8] ), .I1(\preSatVoltage[10] ), 
            .I2(\preSatVoltage[9] ), .I3(n20180), .O(n22));
    defparam i1213_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut_adj_218 (.I0(\preSatVoltage[12] ), .I1(\preSatVoltage[13] ), 
            .I2(n22), .I3(\preSatVoltage[11] ), .O(n19450));
    defparam i1_4_lut_adj_218.LUT_INIT = 16'h8880;
    SB_LUT4 i1_4_lut_adj_219 (.I0(\preSatVoltage[15] ), .I1(\preSatVoltage[16] ), 
            .I2(n19450), .I3(\preSatVoltage[14] ), .O(n19743));
    defparam i1_4_lut_adj_219.LUT_INIT = 16'h8880;
    SB_LUT4 i1_4_lut_adj_220 (.I0(\preSatVoltage[19] ), .I1(\preSatVoltage[18] ), 
            .I2(n19743), .I3(\preSatVoltage[17] ), .O(n20108));
    defparam i1_4_lut_adj_220.LUT_INIT = 16'h8880;
    SB_LUT4 i1_4_lut_adj_221 (.I0(\preSatVoltage[22] ), .I1(n20108), .I2(\preSatVoltage[21] ), 
            .I3(\preSatVoltage[20] ), .O(n20092));
    defparam i1_4_lut_adj_221.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_222 (.I0(\preSatVoltage[25] ), .I1(\preSatVoltage[24] ), 
            .I2(n20092), .I3(\preSatVoltage[23] ), .O(n19914));
    defparam i1_4_lut_adj_222.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_223 (.I0(\preSatVoltage[28] ), .I1(\preSatVoltage[27] ), 
            .I2(\preSatVoltage[26] ), .I3(n19914), .O(n19920));
    defparam i1_4_lut_adj_223.LUT_INIT = 16'hfffe;
    SB_LUT4 i12830_4_lut (.I0(\preSatVoltage[29] ), .I1(\Voltage_1[31] ), 
            .I2(\preSatVoltage[30] ), .I3(n19920), .O(Out_31__N_332));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[37:72])
    defparam i12830_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_224 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[11]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n426));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_224.LUT_INIT = 16'h4440;
    SB_LUT4 i13215_2_lut_3_lut (.I0(\preSatVoltage[22] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[13] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13215_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_225 (.I0(\preSatVoltage[22] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n685));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_225.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_226 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[3]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n402));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_226.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_227 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[12]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n429));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_227.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_228 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[13]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n432));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_228.LUT_INIT = 16'h4440;
    SB_LUT4 i3_4_lut_adj_229 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[8]), .O(n26));
    defparam i3_4_lut_adj_229.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_230 (.I0(\preSatVoltage[16] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n391));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_230.LUT_INIT = 16'h00d0;
    SB_LUT4 i3_4_lut_adj_231 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[7]), .O(n23));
    defparam i3_4_lut_adj_231.LUT_INIT = 16'h0400;
    SB_LUT4 i13209_2_lut_3_lut (.I0(\preSatVoltage[16] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[7] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13209_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_232 (.I0(\preSatVoltage[16] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n391_adj_22));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_232.LUT_INIT = 16'h00d0;
    SB_LUT4 equal_13244_i21_2_lut_3_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(n21));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam equal_13244_i21_2_lut_3_lut.LUT_INIT = 16'h5858;
    SB_LUT4 Q_15__I_0_11_i369_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(\Product_mul_temp[26] ), .O(n576));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_11_i369_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i389_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[12]), .O(n576_adj_23));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i389_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i387_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[11]), .O(n573));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i387_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i385_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[10]), .O(n570));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i385_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i383_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[9]), .O(n567));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i383_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i13214_2_lut_3_lut (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[12] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13214_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 Q_15__I_0_i381_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[8]), .O(n564));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i381_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_233 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[4]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n405));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_233.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_234 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n628));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_234.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_235 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), .O(n625));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_235.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_236 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n622));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_236.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_237 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[14]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n435));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_237.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_238 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), .O(n619));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_238.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_239 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), .O(n616));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_239.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_240 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[8]), .I3(Out_31__N_332), .O(n613));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_240.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_241 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), .O(n610));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_241.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_242 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[6]), .I3(Out_31__N_332), .O(n607));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_242.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_243 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n601));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_243.LUT_INIT = 16'h00e0;
    SB_LUT4 Q_15__I_0_i379_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[7]), .O(n561));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i379_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_244 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n598));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_244.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_245 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n595));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_245.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_246 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n592));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_246.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_247 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n589));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_247.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_248 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n604));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_248.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_249 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), .O(n631));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_249.LUT_INIT = 16'h00e0;
    SB_LUT4 i13210_2_lut_3_lut (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[8] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13210_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 Q_15__I_0_i377_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[6]), .O(n558));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i377_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i3_4_lut_adj_250 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[6]), .O(n20));
    defparam i3_4_lut_adj_250.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_251 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[6]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[14] ), .O(n264));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_251.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_252 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[6]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n117));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_252.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_253 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[6]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n411));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_253.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_254 (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n587));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_254.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_255 (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n587_adj_24));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_255.LUT_INIT = 16'h00d0;
    SB_LUT4 Q_15__I_0_i393_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[14]), .O(n582));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i393_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_256 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[0]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n393));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_256.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_257 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n408));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_257.LUT_INIT = 16'h00e0;
    SB_LUT4 Q_15__I_0_i375_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[5]), .O(n555));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i375_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i373_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[4]), .O(n552));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i373_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i371_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[3]), .O(n549));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i371_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_258 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[1]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n396));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_258.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_259 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[2]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n399));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_259.LUT_INIT = 16'h4440;
    SB_LUT4 Q_15__I_0_i369_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[2]), .O(n546));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i369_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i13216_2_lut_3_lut (.I0(\preSatVoltage[23] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\qVoltage[14] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13216_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 Q_15__I_0_i367_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[1]), .O(n543));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i367_2_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 Q_15__I_0_i365_2_lut_4_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(Look_Up_Table_out1_1[0]), .O(n540));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam Q_15__I_0_i365_2_lut_4_lut.LUT_INIT = 16'hf200;
    
endmodule
//
// Verilog Description of module D_Current_Control_U1
//

module D_Current_Control_U1 (GND_net, \Product_mul_temp[26] , \Error_sub_temp[31] , 
            n146, \preSatVoltage[23] , \preSatVoltage[19] , n794, pin3_clk_16mhz_N_keep, 
            \preSatVoltage[12] , n141, \Error_sub_temp[30] , Out_31__N_333, 
            Out_31__N_332, \dVoltage[5] , \dVoltage[2] , \dVoltage[8] , 
            \dVoltage[12] , \dVoltage[15] , \dVoltage[13] , \dVoltage[6] , 
            \dVoltage[9] , \dVoltage[11] , \dVoltage[10] , \dVoltage[7] , 
            \dVoltage[3] , \dVoltage[14] , \preSatVoltage[10] , n142, 
            n14349, n14348, n14347, n14346, n14345, n14344, n14343, 
            n14342, n14341, n14340, n14339, n14338, n14320, n14337, 
            n14336, n14335, n14334, n14333, n14332, n14331, n14330, 
            n14329, \Add_add_temp[34] , \Add_add_temp[33] , \Add_add_temp[32] , 
            \Add_add_temp[31] , \Add_add_temp[30] , \Add_add_temp[29] , 
            \Add_add_temp[28] , \Add_add_temp[27] , \Add_add_temp[26] , 
            \Add_add_temp[25] , \Add_add_temp[24] , \Add_add_temp[23] , 
            \Add_add_temp[22] , \Add_add_temp[21] , \Add_add_temp[20] , 
            \Add_add_temp[19] , \Add_add_temp[18] , \Add_add_temp[17] , 
            \Add_add_temp[16] , \Add_add_temp[15] , \Add_add_temp[14] , 
            \Add_add_temp[13] , \Add_add_temp[12] , \Add_add_temp[11] , 
            \Add_add_temp[10] , \Add_add_temp[9] , \Add_add_temp[8] , 
            \Add_add_temp[7] , \Add_add_temp[6] , \Add_add_temp[5] , \Add_add_temp[4] , 
            n14328, n14327, n14326, n14322, n793, n14325, n19782, 
            n14324, n31, n14323, n14321, Saturate_out1_31__N_267, 
            Saturate_out1_31__N_266, \dCurrent[3] , \dCurrent[4] , \dCurrent[5] , 
            \dCurrent[6] , \dCurrent[7] , \dCurrent[8] , \dCurrent[9] , 
            \dCurrent[10] , \dCurrent[11] , \dCurrent[12] , \dCurrent[13] , 
            \dCurrent[14] , \dCurrent[15] , \dCurrent[16] , \dCurrent[17] , 
            \dCurrent[18] , \dCurrent[19] , \dCurrent[20] , \dCurrent[21] , 
            \dCurrent[22] , \dCurrent[23] , \dCurrent[24] , \dCurrent[25] , 
            \dCurrent[26] , \dCurrent[27] , \dCurrent[28] , \dCurrent[29] , 
            \dCurrent[30] , \dCurrent[31] , n342, Look_Up_Table_out1_1, 
            n342_adj_10, n114, n408, n14, n604, n685, n685_adj_11, 
            n417, n123, n613, n429, n135, n625, n587, n587_adj_12, 
            n399, n426, n414, n432, n393, n405, n402, n396, 
            n420, n423, n44, n489, n8, n489_adj_13, n20, n126, 
            n616, n391, n391_adj_14, n19576, n129, n619, n11, 
            n35, n19352, n26, \Product3_mul_temp[2] , n120, n111, 
            n102, n99, n108, n138, n132, n105, n610, n595, n23, 
            n622, n41, n601, n592, n598, n589, n628, n32, n538, 
            n29, n17, n71, n83, n59, n50, n92, n68, n62, n53, 
            n65, n38, n56, n80, n244, n233, n200, n203, n86, 
            n77, n197, n239, n206, n86_adj_15, n215, n89, n74, 
            n227, n233_adj_16, n224, n221, n209, n236, n230, n244_adj_17, 
            n212, n218, n279, n270, n267, n255, n285, n264, 
            n258, n249, n246, n273, n282, n261, n19681, n288, 
            n276, n252, n789, n785, n765, n753, n741, n757, 
            n745, n761, n195, n737, n749, n781, n777, n773, 
            n769, n19684, n435, n141_adj_18, n631, n117, n411, 
            n607) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Product_mul_temp[26] ;
    output \Error_sub_temp[31] ;
    output n146;
    output \preSatVoltage[23] ;
    output \preSatVoltage[19] ;
    input n794;
    input pin3_clk_16mhz_N_keep;
    output \preSatVoltage[12] ;
    input n141;
    output \Error_sub_temp[30] ;
    output Out_31__N_333;
    output Out_31__N_332;
    output \dVoltage[5] ;
    output \dVoltage[2] ;
    output \dVoltage[8] ;
    output \dVoltage[12] ;
    output \dVoltage[15] ;
    output \dVoltage[13] ;
    output \dVoltage[6] ;
    output \dVoltage[9] ;
    output \dVoltage[11] ;
    output \dVoltage[10] ;
    output \dVoltage[7] ;
    output \dVoltage[3] ;
    output \dVoltage[14] ;
    output \preSatVoltage[10] ;
    input n142;
    input n14349;
    input n14348;
    input n14347;
    input n14346;
    input n14345;
    input n14344;
    input n14343;
    input n14342;
    input n14341;
    input n14340;
    input n14339;
    input n14338;
    input n14320;
    input n14337;
    input n14336;
    input n14335;
    input n14334;
    input n14333;
    input n14332;
    input n14331;
    input n14330;
    input n14329;
    output \Add_add_temp[34] ;
    output \Add_add_temp[33] ;
    output \Add_add_temp[32] ;
    output \Add_add_temp[31] ;
    output \Add_add_temp[30] ;
    output \Add_add_temp[29] ;
    output \Add_add_temp[28] ;
    output \Add_add_temp[27] ;
    output \Add_add_temp[26] ;
    output \Add_add_temp[25] ;
    output \Add_add_temp[24] ;
    output \Add_add_temp[23] ;
    output \Add_add_temp[22] ;
    output \Add_add_temp[21] ;
    output \Add_add_temp[20] ;
    output \Add_add_temp[19] ;
    output \Add_add_temp[18] ;
    output \Add_add_temp[17] ;
    output \Add_add_temp[16] ;
    output \Add_add_temp[15] ;
    output \Add_add_temp[14] ;
    output \Add_add_temp[13] ;
    output \Add_add_temp[12] ;
    output \Add_add_temp[11] ;
    output \Add_add_temp[10] ;
    output \Add_add_temp[9] ;
    output \Add_add_temp[8] ;
    output \Add_add_temp[7] ;
    output \Add_add_temp[6] ;
    output \Add_add_temp[5] ;
    output \Add_add_temp[4] ;
    input n14328;
    input n14327;
    input n14326;
    input n14322;
    input n793;
    input n14325;
    input n19782;
    input n14324;
    input n31;
    input n14323;
    input n14321;
    output Saturate_out1_31__N_267;
    output Saturate_out1_31__N_266;
    input \dCurrent[3] ;
    input \dCurrent[4] ;
    input \dCurrent[5] ;
    input \dCurrent[6] ;
    input \dCurrent[7] ;
    input \dCurrent[8] ;
    input \dCurrent[9] ;
    input \dCurrent[10] ;
    input \dCurrent[11] ;
    input \dCurrent[12] ;
    input \dCurrent[13] ;
    input \dCurrent[14] ;
    input \dCurrent[15] ;
    input \dCurrent[16] ;
    input \dCurrent[17] ;
    input \dCurrent[18] ;
    input \dCurrent[19] ;
    input \dCurrent[20] ;
    input \dCurrent[21] ;
    input \dCurrent[22] ;
    input \dCurrent[23] ;
    input \dCurrent[24] ;
    input \dCurrent[25] ;
    input \dCurrent[26] ;
    input \dCurrent[27] ;
    input \dCurrent[28] ;
    input \dCurrent[29] ;
    input \dCurrent[30] ;
    input \dCurrent[31] ;
    output n342;
    input [15:0]Look_Up_Table_out1_1;
    output n342_adj_10;
    output n114;
    output n408;
    output n14;
    output n604;
    output n685;
    output n685_adj_11;
    output n417;
    output n123;
    output n613;
    output n429;
    output n135;
    output n625;
    output n587;
    output n587_adj_12;
    output n399;
    output n426;
    output n414;
    output n432;
    output n393;
    output n405;
    output n402;
    output n396;
    output n420;
    output n423;
    output n44;
    output n489;
    output n8;
    output n489_adj_13;
    output n20;
    output n126;
    output n616;
    output n391;
    output n391_adj_14;
    output n19576;
    output n129;
    output n619;
    output n11;
    output n35;
    output n19352;
    output n26;
    output \Product3_mul_temp[2] ;
    output n120;
    output n111;
    output n102;
    output n99;
    output n108;
    output n138;
    output n132;
    output n105;
    output n610;
    output n595;
    output n23;
    output n622;
    output n41;
    output n601;
    output n592;
    output n598;
    output n589;
    output n628;
    output n32;
    output n538;
    output n29;
    output n17;
    output n71;
    output n83;
    output n59;
    output n50;
    output n92;
    output n68;
    output n62;
    output n53;
    output n65;
    output n38;
    output n56;
    output n80;
    output n244;
    output n233;
    output n200;
    output n203;
    output n86;
    output n77;
    output n197;
    output n239;
    output n206;
    output n86_adj_15;
    output n215;
    output n89;
    output n74;
    output n227;
    output n233_adj_16;
    output n224;
    output n221;
    output n209;
    output n236;
    output n230;
    output n244_adj_17;
    output n212;
    output n218;
    output n279;
    output n270;
    output n267;
    output n255;
    output n285;
    output n264;
    output n258;
    output n249;
    output n246;
    output n273;
    output n282;
    output n261;
    output n19681;
    output n288;
    output n276;
    output n252;
    output n789;
    output n785;
    output n765;
    output n753;
    output n741;
    output n757;
    output n745;
    output n761;
    output n195;
    output n737;
    output n749;
    output n781;
    output n777;
    output n773;
    output n769;
    output n19684;
    output n435;
    output n141_adj_18;
    output n631;
    output n117;
    output n411;
    output n607;
    
    
    wire n17581;
    wire [14:0]n837;
    
    wire n111_c, n17582, n17593, n17594;
    wire [31:0]preSatVoltage;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(55[22:35])
    wire [31:0]Proportional_Gain_mul_temp;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(46[22:48])
    wire [31:0]currentControlITerm;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(59[21:40])
    
    wire n15591, n17526;
    wire [14:0]n833;
    
    wire n17527, n17609;
    wire [14:0]n838;
    
    wire n757_c, n759, n17558;
    wire [14:0]n835;
    
    wire n105_c, n17559, n17525, n17617;
    wire [14:0]n839;
    
    wire n117_c, n17618;
    wire [14:0]n834;
    
    wire n17563, n17574;
    wire [14:0]n836;
    
    wire n108_c, n17575, n17524;
    wire [14:0]n840;
    
    wire n120_c, n17635, n17654;
    wire [14:0]n841;
    
    wire n769_c, n771, n17523, n15592, n17522, n17586, n17521, 
        n17592, n114_c, n17608, n17616, n17552, n17553;
    wire [31:0]Switch_out1;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(58[22:33])
    wire [14:0]n844;
    
    wire n783, n17723, Not_Equal_relop1_N_201, n17636, n17623, n123_c, 
        n17653, n17724, n17587, n17624, n17652, n17899, n17900, 
        n15590;
    wire [14:0]n835_adj_564;
    wire [14:0]n836_adj_565;
    
    wire n138_c, n17777, n17778, n135_c, n17776, n15589, n15588, 
        n15587, n15586, n15585, n15584, n102_c;
    wire [14:0]n843;
    
    wire n779, n17722, n17585, n17541, n796, n17520, n17634, n17651, 
        n791, n17519, n15583, n17545, n17546, n17557;
    wire [31:0]Saturate_out1;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(64[22:35])
    wire [14:0]n842;
    
    wire n775, n17721, n132_c, n17775;
    wire [14:0]n845;
    
    wire n787, n17518;
    wire [14:0]n844_adj_566;
    
    wire n783_adj_349, n17517, n129_c, n17774;
    wire [14:0]n843_adj_567;
    
    wire n779_adj_352, n17516, n17607, n17615;
    wire [14:0]n841_adj_568;
    
    wire n771_adj_353, n17720, n17622;
    wire [14:0]n840_adj_569;
    
    wire n767, n17719, n17650;
    wire [14:0]n839_adj_570;
    
    wire n763, n17718;
    wire [14:0]n838_adj_571;
    
    wire n759_adj_354, n17717;
    wire [14:0]n837_adj_572;
    
    wire n755, n17716, n17633, n17606, n17591, n17554, n15582, 
        n15581, n17547, n17564, n17573, n15580;
    wire [14:0]n842_adj_573;
    
    wire n775_adj_357, n17515, n15579, n15578, n15577, n17548, n17806, 
        n17807;
    wire [32:0]Error_sub_temp;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(44[22:36])
    
    wire n4, n17808;
    wire [14:0]n834_adj_574;
    
    wire n17739, n126_c, n17773, n17742, n17743, n17740, n17741, 
        n20546, n20550, n20548, n20556, n15, n20554, n20560, n20562, 
        n20568, n20566, n751, n17715, n785_c, n20574, n14_c, n20576, 
        n20572, n19727, n20198, n19858, n17649, n17772, n15576, 
        n12, n19269, n15575, n15574, n20196, n15573, n20194, n15572, 
        n20192, n15571, n20190, n15570, n20188, n15569, n20186, 
        n15568, n20184;
    wire [31:0]Voltage_1;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(56[22:31])
    
    wire n15597, n15593, n777_c, n17275, n17274, n17273, n17756, 
        n17757, n17272, n17271, n17270, n789_c, n17269, n17268, 
        n17267, n17266, n16003, n16002, n16001, n16000, n15999, 
        n15998, n15997, n15996, n15995, n15994, n15993, n15992, 
        n15991, n15990, n15989, n15988, n15987, n15986, n15985, 
        n15984, n15983, n15982, n15981, n15980, n15979, n15978, 
        n15977, n15976, n15975, n15974, n17771, n19273, n17738, 
        n17770, n17805, n17824, n747, n17714, n17823, n17737, 
        n743, n17713, n17769;
    wire [14:0]n833_adj_575;
    
    wire n8265, n17712, n17804, n17822, n17768, n17514, n15973, 
        n17753, n17803, n17562, n17898, n17821, n17802, n17767, 
        n767_adj_382, n17513, n17766, n763_adj_386, n17512, n17901, 
        n17897, n17572, n17895, n17571, n17570, n17894, n17569, 
        n17568, n17549, n17556, n18172, n18171, n18170, n18169, 
        n18168, n18167, n17801, n17511, n755_adj_404, n17510, n751_adj_406, 
        n17509, n747_adj_408, n17508, n743_adj_410, n17507, n739, 
        n17506, n17505;
    wire [14:0]n832;
    
    wire n17820, n17736, n781_c, n18142, n18141, n18140, n18139, 
        n18138, n18137, n18136, n18135, n773_c, n18133, n18132, 
        n18131, n18130, n18129, n18128, n18127, n18126, n18125, 
        n18124, n18123, n18122;
    wire [14:0]n846;
    
    wire n17955, n795, n17954, n17953, n17952, n17951, n17950, 
        n17949, n765_c, n17948, n761_c, n17947, n17946, n753_c, 
        n17945, n749_c, n17944, n745_c, n17943, n741_c, n17942, 
        n737_c;
    wire [14:0]n845_adj_576;
    
    wire n17940, n791_adj_416, n17939, n17938, n17937, n17936, n17935, 
        n17934, n17933, n17932, n17931, n17930, n17929, n17928, 
        n17927, n17925, n787_adj_421, n17924, n17923, n17922, n17919, 
        n17920, n17921, n17893, n17579, n17892, n17754, n17800, 
        n17711, n17819;
    wire [14:0]n832_adj_577;
    
    wire n17799, n17764, n17818, n17817, n17798, n17752, n17797, 
        n17891, n17751, n17763, n17816, n17762, n17890, n17796, 
        n17889, n17761, n17888, n17815, n17887, n17814, n17542, 
        n17555, n17561, n17567, n17886, n17813, n17578, n17584, 
        n17590, n17621, n17885, n17812, n17632, n17648, n17794, 
        n17811, n17884, n17883, n17882, n17760, n17793, n17809, 
        n17605, n17880, n17879, n17878, n17877, n17876, n17875, 
        n17874, n17540, n17566, n17873, n17577, n17583, n17589, 
        n17759, n17604, n17614, n17872, n17792, n17871, n17631, 
        n17647, n17870, n17791, n17869, n17868, n17867, n15594, 
        n15595, n15596, n17539, n17551, n17560, n17603, n17602, 
        n17601, n17600, n17599, n17598, n17597, n17596, n17646, 
        n17630, n17613, n17790, n17620, n17544, n17749, n17645, 
        n17758, n17789, n17629, n17619, n17854, n17853, n17852, 
        n17628, n17851, n17850, n17849, n17848, n17847, n17846, 
        n17576, n17845, n17538, n17543, n17644, n17844, n17588, 
        n17788, n17612, n17843, n17627, n17643, n17842, n17841, 
        n17748, n17787, n17839, n17642, n17838, n17837, n17836, 
        n17835, n17834, n17833, n17832, n17831, n17786, n17611, 
        n17830, n17537, n17829, n17828, n17785, n17626, n17827, 
        n17826, n17641, n17784, n17747, n17783, n17746, n17755, 
        n17745, n17744, n17782, n17726, n17781, n17725, n17639, 
        n17918, n17638, n17779, n17917, n17637, n17536, n17916, 
        n17915, n17914;
    wire [31:0]n1;
    
    wire n15804, n15803, n15802, n17913, n15801, n15800, n15799, 
        n15798, n15797, n15796, n15795, n17912, n15794, n15793, 
        n15792, n15791, n15790, n15789, n15788, n15787, n15786, 
        n15785, n15784, n15783, n15782, n15781, n17910, n15780, 
        n15779, n15778, n15777, n15776, n15775, VCC_net, n17909, 
        n17908, n17907, n17906, n17905, n17904, n17903, n17902, 
        n20712, n17534, n17533, n17532, n17531, n17530, n17529, 
        n19777, n17528, n20700, n15205, n20670, n19746, n20656, 
        n20648, n20634, n15264, n19723, n20708, n22_adj_519, n20688, 
        n19842, n20666, n20658, n20644, n58;
    
    SB_CARRY paramCurrentControlP_15__I_0_add_565_3 (.CI(n17581), .I0(n837[0]), 
            .I1(n111_c), .CO(n17582));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_15 (.CI(n17593), .I0(n837[12]), 
            .I1(n111_c), .CO(n17594));
    SB_LUT4 add_547_26_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[24]), 
            .I2(currentControlITerm[31]), .I3(n15591), .O(preSatVoltage[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_8 (.CI(n17526), .I0(n833[5]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17527));
    SB_CARRY paramCurrentControlP_15__I_0_add_566_16 (.CI(n17609), .I0(n838[13]), 
            .I1(n757_c), .CO(n759));
    SB_CARRY paramCurrentControlP_15__I_0_add_563_10 (.CI(n17558), .I0(n835[7]), 
            .I1(n105_c), .CO(n17559));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_7_lut (.I0(GND_net), .I1(n833[4]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17525), .O(Proportional_Gain_mul_temp[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_9 (.CI(n17617), .I0(n839[6]), 
            .I1(n117_c), .CO(n17618));
    SB_CARRY paramCurrentControlP_15__I_0_add_561_7 (.CI(n17525), .I0(n833[4]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17526));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_15_lut (.I0(GND_net), .I1(n835[12]), 
            .I2(n105_c), .I3(n17563), .O(n834[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_11 (.CI(n17574), .I0(n836[8]), 
            .I1(n108_c), .CO(n17575));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_6_lut (.I0(GND_net), .I1(n833[3]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17524), .O(Proportional_Gain_mul_temp[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_12_lut (.I0(GND_net), .I1(n840[9]), 
            .I2(n120_c), .I3(n17635), .O(n839[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_6 (.CI(n17524), .I0(n833[3]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17525));
    SB_CARRY paramCurrentControlP_15__I_0_add_569_16 (.CI(n17654), .I0(n841[11]), 
            .I1(n769_c), .CO(n771));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_5_lut (.I0(GND_net), .I1(n833[2]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17523), .O(Proportional_Gain_mul_temp[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_26 (.CI(n15591), .I0(Proportional_Gain_mul_temp[24]), 
            .I1(currentControlITerm[31]), .CO(n15592));
    SB_CARRY paramCurrentControlP_15__I_0_add_561_5 (.CI(n17523), .I0(n833[2]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17524));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_4_lut (.I0(GND_net), .I1(n833[1]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17522), .O(Proportional_Gain_mul_temp[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_4 (.CI(n17522), .I0(n833[1]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17523));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_8_lut (.I0(GND_net), .I1(n837[5]), 
            .I2(n111_c), .I3(n17586), .O(n836[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_3_lut (.I0(GND_net), .I1(n833[0]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17521), .O(Proportional_Gain_mul_temp[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_14_lut (.I0(GND_net), .I1(n837[11]), 
            .I2(n111_c), .I3(n17592), .O(n836[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_15_lut (.I0(GND_net), .I1(n838[12]), 
            .I2(n114_c), .I3(n17608), .O(n837[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_i66_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(\Error_sub_temp[31] ), .I2(GND_net), .I3(GND_net), .O(n146));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i66_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_8_lut (.I0(GND_net), .I1(n839[5]), 
            .I2(n117_c), .I3(n17616), .O(n838[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_4 (.CI(n17552), .I0(n835[1]), 
            .I1(n105_c), .CO(n17553));
    SB_LUT4 add_4257_14_lut (.I0(Not_Equal_relop1_N_201), .I1(n844[14]), 
            .I2(n783), .I3(n17723), .O(Switch_out1[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_12 (.CI(n17635), .I0(n840[9]), 
            .I1(n120_c), .CO(n17636));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_15_lut (.I0(GND_net), .I1(n839[12]), 
            .I2(n117_c), .I3(n17623), .O(n838[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_15 (.CI(n17608), .I0(n838[12]), 
            .I1(n114_c), .CO(n17609));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_15_lut (.I0(GND_net), .I1(n841[11]), 
            .I2(n123_c), .I3(n17653), .O(n840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_15 (.CI(n17653), .I0(n841[11]), 
            .I1(n123_c), .CO(n17654));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_8 (.CI(n17616), .I0(n839[5]), 
            .I1(n117_c), .CO(n17617));
    SB_CARRY add_4257_14 (.CI(n17723), .I0(n844[14]), .I1(n783), .CO(n17724));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_8 (.CI(n17586), .I0(n837[5]), 
            .I1(n111_c), .CO(n17587));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_15 (.CI(n17623), .I0(n839[12]), 
            .I1(n117_c), .CO(n17624));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_14_lut (.I0(GND_net), .I1(n841[11]), 
            .I2(n123_c), .I3(n17652), .O(n840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_14 (.CI(n17652), .I0(n841[11]), 
            .I1(n123_c), .CO(n17653));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_2_lut (.I0(GND_net), .I1(n114_c), 
            .I2(n111_c), .I3(GND_net), .O(n836[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_5 (.CI(n17899), .I0(n844[2]), 
            .I1(n111_c), .CO(n17900));
    SB_LUT4 add_547_25_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[23]), 
            .I2(currentControlITerm[31]), .I3(n15590), .O(preSatVoltage[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_564_14_lut (.I0(GND_net), .I1(n836_adj_565[11]), 
            .I2(n138_c), .I3(n17777), .O(n835_adj_564[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_14 (.CI(n17777), .I0(n836_adj_565[11]), 
            .I1(n138_c), .CO(n17778));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_13_lut (.I0(GND_net), .I1(n836_adj_565[10]), 
            .I2(n135_c), .I3(n17776), .O(n835_adj_564[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_3 (.CI(n17521), .I0(n833[0]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17522));
    SB_CARRY add_547_25 (.CI(n15590), .I0(Proportional_Gain_mul_temp[23]), 
            .I1(currentControlITerm[31]), .CO(n15591));
    SB_LUT4 add_547_24_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[22]), 
            .I2(currentControlITerm[30]), .I3(n15589), .O(\preSatVoltage[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_24 (.CI(n15589), .I0(Proportional_Gain_mul_temp[22]), 
            .I1(currentControlITerm[30]), .CO(n15590));
    SB_LUT4 add_547_23_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[21]), 
            .I2(currentControlITerm[29]), .I3(n15588), .O(preSatVoltage[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_23 (.CI(n15588), .I0(Proportional_Gain_mul_temp[21]), 
            .I1(currentControlITerm[29]), .CO(n15589));
    SB_LUT4 add_547_22_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[20]), 
            .I2(currentControlITerm[28]), .I3(n15587), .O(preSatVoltage[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_22 (.CI(n15587), .I0(Proportional_Gain_mul_temp[20]), 
            .I1(currentControlITerm[28]), .CO(n15588));
    SB_LUT4 add_547_21_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[19]), 
            .I2(currentControlITerm[27]), .I3(n15586), .O(preSatVoltage[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_21 (.CI(n15586), .I0(Proportional_Gain_mul_temp[19]), 
            .I1(currentControlITerm[27]), .CO(n15587));
    SB_LUT4 add_547_20_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[18]), 
            .I2(currentControlITerm[26]), .I3(n15585), .O(\preSatVoltage[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_20 (.CI(n15585), .I0(Proportional_Gain_mul_temp[18]), 
            .I1(currentControlITerm[26]), .CO(n15586));
    SB_LUT4 add_547_19_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[17]), 
            .I2(currentControlITerm[25]), .I3(n15584), .O(preSatVoltage[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_19 (.CI(n15584), .I0(Proportional_Gain_mul_temp[17]), 
            .I1(currentControlITerm[25]), .CO(n15585));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_2_lut (.I0(GND_net), .I1(n102_c), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(GND_net), .O(Proportional_Gain_mul_temp[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_2 (.CI(GND_net), .I0(n102_c), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17521));
    SB_LUT4 add_4257_13_lut (.I0(Not_Equal_relop1_N_201), .I1(n843[14]), 
            .I2(n779), .I3(n17722), .O(Switch_out1[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_7_lut (.I0(GND_net), .I1(n837[4]), 
            .I2(n111_c), .I3(n17585), .O(n836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_8_lut (.I0(GND_net), .I1(n834[5]), 
            .I2(n102_c), .I3(n17541), .O(n833[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_17_lut (.I0(GND_net), .I1(n796), .I2(GND_net), .I3(n17520), 
            .O(Proportional_Gain_mul_temp[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_11_lut (.I0(GND_net), .I1(n840[8]), 
            .I2(n120_c), .I3(n17634), .O(n839[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_13_lut (.I0(GND_net), .I1(n841[10]), 
            .I2(n123_c), .I3(n17651), .O(n840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_16_lut (.I0(GND_net), .I1(n794), .I2(n791), .I3(n17519), 
            .O(Proportional_Gain_mul_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_547_18_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[16]), 
            .I2(currentControlITerm[24]), .I3(n15583), .O(preSatVoltage[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_18 (.CI(n15583), .I0(Proportional_Gain_mul_temp[16]), 
            .I1(currentControlITerm[24]), .CO(n15584));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_4_lut (.I0(GND_net), .I1(n835[1]), 
            .I2(n105_c), .I3(n17552), .O(n834[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_14 (.CI(n17592), .I0(n837[11]), 
            .I1(n111_c), .CO(n17593));
    SB_CARRY paramCurrentControlP_15__I_0_add_562_12 (.CI(n17545), .I0(n834[9]), 
            .I1(n102_c), .CO(n17546));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_9_lut (.I0(GND_net), .I1(n835[6]), 
            .I2(n105_c), .I3(n17557), .O(n834[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4257_13 (.CI(n17722), .I0(n843[14]), .I1(n779), .CO(n17723));
    SB_DFF currentControlITerm_i31 (.Q(currentControlITerm[31]), .C(pin3_clk_16mhz_N_keep), 
           .D(Saturate_out1[31]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_CARRY Error_sub_temp_31__I_0_add_564_13 (.CI(n17776), .I0(n836_adj_565[10]), 
            .I1(n135_c), .CO(n17777));
    SB_LUT4 add_4257_12_lut (.I0(Not_Equal_relop1_N_201), .I1(n842[14]), 
            .I2(n775), .I3(n17721), .O(Switch_out1[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4257_12 (.CI(n17721), .I0(n842[14]), .I1(n775), .CO(n17722));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_12_lut (.I0(GND_net), .I1(n836_adj_565[9]), 
            .I2(n132_c), .I3(n17775), .O(n835_adj_564[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_12 (.CI(n17775), .I0(n836_adj_565[9]), 
            .I1(n132_c), .CO(n17776));
    SB_CARRY add_3099_16 (.CI(n17519), .I0(n794), .I1(n791), .CO(n17520));
    SB_LUT4 add_3099_15_lut (.I0(GND_net), .I1(n845[14]), .I2(n787), .I3(n17518), 
            .O(Proportional_Gain_mul_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_15 (.CI(n17518), .I0(n845[14]), .I1(n787), .CO(n17519));
    SB_LUT4 add_3099_14_lut (.I0(GND_net), .I1(n844_adj_566[14]), .I2(n783_adj_349), 
            .I3(n17517), .O(Proportional_Gain_mul_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_14 (.CI(n17517), .I0(n844_adj_566[14]), .I1(n783_adj_349), 
            .CO(n17518));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_11_lut (.I0(GND_net), .I1(n836_adj_565[8]), 
            .I2(n129_c), .I3(n17774), .O(n835_adj_564[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_13_lut (.I0(GND_net), .I1(n843_adj_567[14]), .I2(n779_adj_352), 
            .I3(n17516), .O(Proportional_Gain_mul_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_13 (.CI(n17516), .I0(n843_adj_567[14]), .I1(n779_adj_352), 
            .CO(n17517));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_14_lut (.I0(GND_net), .I1(n838[11]), 
            .I2(n114_c), .I3(n17607), .O(n837[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_13 (.CI(n17651), .I0(n841[10]), 
            .I1(n123_c), .CO(n17652));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_7_lut (.I0(GND_net), .I1(n839[4]), 
            .I2(n117_c), .I3(n17615), .O(n838[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4257_11_lut (.I0(Not_Equal_relop1_N_201), .I1(n841_adj_568[14]), 
            .I2(n771_adj_353), .I3(n17720), .O(Switch_out1[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_14_lut (.I0(GND_net), .I1(n839[11]), 
            .I2(n117_c), .I3(n17622), .O(n838[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4257_11 (.CI(n17720), .I0(n841_adj_568[14]), .I1(n771_adj_353), 
            .CO(n17721));
    SB_LUT4 add_4257_10_lut (.I0(Not_Equal_relop1_N_201), .I1(n840_adj_569[14]), 
            .I2(n767), .I3(n17719), .O(Switch_out1[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4257_10 (.CI(n17719), .I0(n840_adj_569[14]), .I1(n767), 
            .CO(n17720));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_12_lut (.I0(GND_net), .I1(n841[9]), 
            .I2(n123_c), .I3(n17650), .O(n840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4257_9_lut (.I0(Not_Equal_relop1_N_201), .I1(n839_adj_570[14]), 
            .I2(n763), .I3(n17718), .O(Switch_out1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_11 (.CI(n17634), .I0(n840[8]), 
            .I1(n120_c), .CO(n17635));
    SB_CARRY add_4257_9 (.CI(n17718), .I0(n839_adj_570[14]), .I1(n763), 
            .CO(n17719));
    SB_LUT4 add_4257_8_lut (.I0(Not_Equal_relop1_N_201), .I1(n838_adj_571[14]), 
            .I2(n759_adj_354), .I3(n17717), .O(Switch_out1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_12 (.CI(n17650), .I0(n841[9]), 
            .I1(n123_c), .CO(n17651));
    SB_CARRY add_4257_8 (.CI(n17717), .I0(n838_adj_571[14]), .I1(n759_adj_354), 
            .CO(n17718));
    SB_LUT4 add_4257_7_lut (.I0(Not_Equal_relop1_N_201), .I1(n837_adj_572[14]), 
            .I2(n755), .I3(n17716), .O(Switch_out1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_12_lut (.I0(GND_net), .I1(n834[9]), 
            .I2(n102_c), .I3(n17545), .O(n833[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_10_lut (.I0(GND_net), .I1(n840[7]), 
            .I2(n120_c), .I3(n17633), .O(n839[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_14 (.CI(n17607), .I0(n838[11]), 
            .I1(n114_c), .CO(n17608));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_13_lut (.I0(GND_net), .I1(n838[10]), 
            .I2(n114_c), .I3(n17606), .O(n837[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_10 (.CI(n17633), .I0(n840[7]), 
            .I1(n120_c), .CO(n17634));
    SB_CARRY add_4257_7 (.CI(n17716), .I0(n837_adj_572[14]), .I1(n755), 
            .CO(n17717));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_2 (.CI(GND_net), .I0(n114_c), 
            .I1(n111_c), .CO(n17581));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_13_lut (.I0(GND_net), .I1(n837[10]), 
            .I2(n111_c), .I3(n17591), .O(n836[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_5 (.CI(n17553), .I0(n835[2]), 
            .I1(n105_c), .CO(n17554));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_5_lut (.I0(GND_net), .I1(n835[2]), 
            .I2(n105_c), .I3(n17553), .O(n834[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_547_17_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[15]), 
            .I2(currentControlITerm[23]), .I3(n15582), .O(preSatVoltage[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_17 (.CI(n15582), .I0(Proportional_Gain_mul_temp[15]), 
            .I1(currentControlITerm[23]), .CO(n15583));
    SB_LUT4 add_547_16_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[14]), 
            .I2(currentControlITerm[22]), .I3(n15581), .O(preSatVoltage[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_16 (.CI(n15581), .I0(Proportional_Gain_mul_temp[14]), 
            .I1(currentControlITerm[22]), .CO(n15582));
    SB_CARRY paramCurrentControlP_15__I_0_add_562_13 (.CI(n17546), .I0(n834[10]), 
            .I1(n102_c), .CO(n17547));
    SB_CARRY paramCurrentControlP_15__I_0_add_563_15 (.CI(n17563), .I0(n835[12]), 
            .I1(n105_c), .CO(n17564));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_10_lut (.I0(GND_net), .I1(n836[7]), 
            .I2(n108_c), .I3(n17573), .O(n835[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_547_15_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[13]), 
            .I2(currentControlITerm[21]), .I3(n15580), .O(preSatVoltage[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_12_lut (.I0(GND_net), .I1(n842_adj_573[14]), .I2(n775_adj_357), 
            .I3(n17515), .O(Proportional_Gain_mul_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_15 (.CI(n15580), .I0(Proportional_Gain_mul_temp[13]), 
            .I1(currentControlITerm[21]), .CO(n15581));
    SB_LUT4 add_547_14_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[12]), 
            .I2(currentControlITerm[20]), .I3(n15579), .O(preSatVoltage[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_14 (.CI(n15579), .I0(Proportional_Gain_mul_temp[12]), 
            .I1(currentControlITerm[20]), .CO(n15580));
    SB_LUT4 add_547_13_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[11]), 
            .I2(currentControlITerm[19]), .I3(n15578), .O(\preSatVoltage[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_13 (.CI(n15578), .I0(Proportional_Gain_mul_temp[11]), 
            .I1(currentControlITerm[19]), .CO(n15579));
    SB_LUT4 add_547_12_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[10]), 
            .I2(currentControlITerm[18]), .I3(n15577), .O(preSatVoltage[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_13_lut (.I0(GND_net), .I1(n834[10]), 
            .I2(n102_c), .I3(n17546), .O(n833[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_14 (.CI(n17547), .I0(n834[11]), 
            .I1(n102_c), .CO(n17548));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_14_lut (.I0(GND_net), .I1(n834[11]), 
            .I2(n102_c), .I3(n17547), .O(n833[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_13 (.CI(n17806), .I0(n838_adj_571[10]), 
            .I1(n135_c), .CO(n17807));
    SB_LUT4 i11961_4_lut (.I0(Error_sub_temp[29]), .I1(n138_c), .I2(n141), 
            .I3(\Error_sub_temp[30] ), .O(n4));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i11961_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 Error_sub_temp_31__I_0_add_566_15_lut (.I0(GND_net), .I1(n838_adj_571[12]), 
            .I2(n141), .I3(n17808), .O(n837_adj_572[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_11 (.CI(n17774), .I0(n836_adj_565[8]), 
            .I1(n129_c), .CO(n17775));
    SB_LUT4 paramCurrentControlP_15__I_0_i51_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[24]), .I2(GND_net), .I3(GND_net), .O(n123_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Error_sub_temp_31__I_0_add_562_6_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[3]), .I2(n114_c), .I3(n17739), .O(Switch_out1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Error_sub_temp_31__I_0_add_564_10_lut (.I0(GND_net), .I1(n836_adj_565[7]), 
            .I2(n126_c), .I3(n17773), .O(n835_adj_564[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_9 (.CI(n17742), .I0(n834_adj_574[6]), 
            .I1(n123_c), .CO(n17743));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_7_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[4]), .I2(n117_c), .I3(n17740), .O(Switch_out1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11954_3_lut (.I0(\Product_mul_temp[26] ), .I1(\Error_sub_temp[30] ), 
            .I2(Error_sub_temp[29]), .I3(GND_net), .O(n845[0]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i11954_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i2_4_lut (.I0(n141), .I1(n138_c), .I2(Error_sub_temp[29]), 
            .I3(n146), .O(n845[1]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_4_lut.LUT_INIT = 16'h39c6;
    SB_LUT4 Error_sub_temp_31__I_0_add_562_8_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[5]), .I2(n120_c), .I3(n17741), .O(Switch_out1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut (.I0(preSatVoltage[26]), .I1(preSatVoltage[27]), .I2(Out_31__N_333), 
            .I3(Out_31__N_332), .O(n20546));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut.LUT_INIT = 16'hee70;
    SB_LUT4 i1_4_lut_adj_117 (.I0(preSatVoltage[30]), .I1(preSatVoltage[29]), 
            .I2(Out_31__N_333), .I3(Out_31__N_332), .O(n20550));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_117.LUT_INIT = 16'hee70;
    SB_LUT4 i1_4_lut_adj_118 (.I0(preSatVoltage[25]), .I1(preSatVoltage[28]), 
            .I2(Out_31__N_333), .I3(Out_31__N_332), .O(n20548));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_118.LUT_INIT = 16'hee70;
    SB_LUT4 i1_2_lut (.I0(n20550), .I1(n20546), .I2(GND_net), .I3(GND_net), 
            .O(n20556));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_13243_i15_2_lut (.I0(preSatVoltage[14]), .I1(\dVoltage[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam equal_13243_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_119 (.I0(preSatVoltage[11]), .I1(preSatVoltage[17]), 
            .I2(\dVoltage[2] ), .I3(\dVoltage[8] ), .O(n20554));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_119.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_120 (.I0(preSatVoltage[21]), .I1(n20554), .I2(n15), 
            .I3(\dVoltage[12] ), .O(n20560));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_120.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_4_lut_adj_121 (.I0(preSatVoltage[24]), .I1(n20556), .I2(n20548), 
            .I3(\dVoltage[15] ), .O(n20562));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_121.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_4_lut_adj_122 (.I0(preSatVoltage[22]), .I1(preSatVoltage[15]), 
            .I2(\dVoltage[13] ), .I3(\dVoltage[6] ), .O(n20568));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_122.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_123 (.I0(preSatVoltage[18]), .I1(preSatVoltage[20]), 
            .I2(\dVoltage[9] ), .I3(\dVoltage[11] ), .O(n20566));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_123.LUT_INIT = 16'h7bde;
    SB_LUT4 add_4257_6_lut (.I0(Not_Equal_relop1_N_201), .I1(n836_adj_565[14]), 
            .I2(n751), .I3(n17715), .O(Switch_out1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 paramCurrentControlP_15__I_0_i534_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[28]), .I2(GND_net), .I3(GND_net), .O(n785_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i534_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_124 (.I0(n20562), .I1(\preSatVoltage[19] ), .I2(n20560), 
            .I3(\dVoltage[10] ), .O(n20574));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_124.LUT_INIT = 16'hfbfe;
    SB_LUT4 i1_4_lut_adj_125 (.I0(preSatVoltage[16]), .I1(n20568), .I2(n14_c), 
            .I3(\dVoltage[7] ), .O(n20576));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_125.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_4_lut_adj_126 (.I0(\preSatVoltage[12] ), .I1(\preSatVoltage[23] ), 
            .I2(\dVoltage[3] ), .I3(\dVoltage[14] ), .O(n20572));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_126.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_127 (.I0(n20572), .I1(n20576), .I2(n20574), .I3(n20566), 
            .O(n19727));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam i1_4_lut_adj_127.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(\preSatVoltage[10] ), .I1(preSatVoltage[9]), .I2(n20198), 
            .I3(GND_net), .O(n19858));
    defparam i1_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_11_lut (.I0(GND_net), .I1(n841[8]), 
            .I2(n123_c), .I3(n17649), .O(n840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 equal_13243_i62_4_lut (.I0(n19858), .I1(n19727), .I2(Out_31__N_333), 
            .I3(Out_31__N_332), .O(Not_Equal_relop1_N_201));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(105[29:55])
    defparam equal_13243_i62_4_lut.LUT_INIT = 16'h2223;
    SB_CARRY Error_sub_temp_31__I_0_add_564_10 (.CI(n17773), .I0(n836_adj_565[7]), 
            .I1(n126_c), .CO(n17774));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_9_lut (.I0(GND_net), .I1(n836_adj_565[6]), 
            .I2(n123_c), .I3(n17772), .O(n835_adj_564[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_12 (.CI(n15577), .I0(Proportional_Gain_mul_temp[10]), 
            .I1(currentControlITerm[18]), .CO(n15578));
    SB_LUT4 add_547_11_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[9]), 
            .I2(currentControlITerm[17]), .I3(n15576), .O(\preSatVoltage[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_3_lut_3_lut (.I0(n138_c), .I1(n142), .I2(n12), .I3(n12), 
            .O(n19269));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_3_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_CARRY add_547_11 (.CI(n15576), .I0(Proportional_Gain_mul_temp[9]), 
            .I1(currentControlITerm[17]), .CO(n15577));
    SB_LUT4 add_547_10_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[8]), 
            .I2(currentControlITerm[16]), .I3(n15575), .O(preSatVoltage[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_10 (.CI(n15575), .I0(Proportional_Gain_mul_temp[8]), 
            .I1(currentControlITerm[16]), .CO(n15576));
    SB_DFF currentControlITerm_i30 (.Q(currentControlITerm[30]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14349));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 add_547_9_lut (.I0(n20196), .I1(Proportional_Gain_mul_temp[7]), 
            .I2(currentControlITerm[15]), .I3(n15574), .O(n20198)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_9 (.CI(n15574), .I0(Proportional_Gain_mul_temp[7]), 
            .I1(currentControlITerm[15]), .CO(n15575));
    SB_LUT4 add_547_8_lut (.I0(n20194), .I1(Proportional_Gain_mul_temp[6]), 
            .I2(currentControlITerm[14]), .I3(n15573), .O(n20196)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_8 (.CI(n15573), .I0(Proportional_Gain_mul_temp[6]), 
            .I1(currentControlITerm[14]), .CO(n15574));
    SB_LUT4 add_547_7_lut (.I0(n20192), .I1(Proportional_Gain_mul_temp[5]), 
            .I2(currentControlITerm[13]), .I3(n15572), .O(n20194)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_7 (.CI(n15572), .I0(Proportional_Gain_mul_temp[5]), 
            .I1(currentControlITerm[13]), .CO(n15573));
    SB_LUT4 add_547_6_lut (.I0(n20190), .I1(Proportional_Gain_mul_temp[4]), 
            .I2(currentControlITerm[12]), .I3(n15571), .O(n20192)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_6 (.CI(n15571), .I0(Proportional_Gain_mul_temp[4]), 
            .I1(currentControlITerm[12]), .CO(n15572));
    SB_LUT4 add_547_5_lut (.I0(n20188), .I1(Proportional_Gain_mul_temp[3]), 
            .I2(currentControlITerm[11]), .I3(n15570), .O(n20190)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_5 (.CI(n15570), .I0(Proportional_Gain_mul_temp[3]), 
            .I1(currentControlITerm[11]), .CO(n15571));
    SB_LUT4 add_547_4_lut (.I0(n20186), .I1(Proportional_Gain_mul_temp[2]), 
            .I2(currentControlITerm[10]), .I3(n15569), .O(n20188)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_4 (.CI(n15569), .I0(Proportional_Gain_mul_temp[2]), 
            .I1(currentControlITerm[10]), .CO(n15570));
    SB_LUT4 add_547_3_lut (.I0(n20184), .I1(Proportional_Gain_mul_temp[1]), 
            .I2(currentControlITerm[9]), .I3(n15568), .O(n20186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_3 (.CI(n15568), .I0(Proportional_Gain_mul_temp[1]), 
            .I1(currentControlITerm[9]), .CO(n15569));
    SB_LUT4 add_547_2_lut (.I0(preSatVoltage[0]), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(currentControlITerm[8]), .I3(GND_net), .O(n20184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_547_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(currentControlITerm[8]), .CO(n15568));
    SB_DFF currentControlITerm_i29 (.Q(currentControlITerm[29]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14348));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i28 (.Q(currentControlITerm[28]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14347));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i27 (.Q(currentControlITerm[27]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14346));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i26 (.Q(currentControlITerm[26]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14345));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i25 (.Q(currentControlITerm[25]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14344));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i24 (.Q(currentControlITerm[24]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14343));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i23 (.Q(currentControlITerm[23]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14342));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i22 (.Q(currentControlITerm[22]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14341));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i21 (.Q(currentControlITerm[21]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14340));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i20 (.Q(currentControlITerm[20]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14339));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i19 (.Q(currentControlITerm[19]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14338));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i1 (.Q(currentControlITerm[1]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14320));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i18 (.Q(currentControlITerm[18]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14337));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i17 (.Q(currentControlITerm[17]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14336));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i16 (.Q(currentControlITerm[16]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14335));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i15 (.Q(currentControlITerm[15]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14334));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i14 (.Q(currentControlITerm[14]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14333));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i13 (.Q(currentControlITerm[13]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14332));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i12 (.Q(currentControlITerm[12]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14331));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i11 (.Q(currentControlITerm[11]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14330));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 add_547_32_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[30]), 
            .I2(currentControlITerm[31]), .I3(n15597), .O(Voltage_1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_27 (.CI(n15592), .I0(Proportional_Gain_mul_temp[25]), 
            .I1(currentControlITerm[31]), .CO(n15593));
    SB_DFF currentControlITerm_i10 (.Q(currentControlITerm[10]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14329));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_12_lut (.I0(GND_net), .I1(n843_adj_567[7]), 
            .I2(n777_c), .I3(n17275), .O(n842_adj_573[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_12 (.CI(n17275), .I0(n843_adj_567[7]), 
            .I1(n777_c), .CO(n779_adj_352));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_11_lut (.I0(GND_net), .I1(n843_adj_567[7]), 
            .I2(n129_c), .I3(n17274), .O(n842_adj_573[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_11 (.CI(n17274), .I0(n843_adj_567[7]), 
            .I1(n129_c), .CO(n17275));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_10_lut (.I0(GND_net), .I1(n843_adj_567[7]), 
            .I2(n129_c), .I3(n17273), .O(n842_adj_573[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_8 (.CI(n17756), .I0(n835_adj_564[5]), 
            .I1(n120_c), .CO(n17757));
    SB_CARRY paramCurrentControlP_15__I_0_add_571_10 (.CI(n17273), .I0(n843_adj_567[7]), 
            .I1(n129_c), .CO(n17274));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_9_lut (.I0(GND_net), .I1(n843_adj_567[6]), 
            .I2(n129_c), .I3(n17272), .O(n842_adj_573[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_9 (.CI(n17272), .I0(n843_adj_567[6]), 
            .I1(n129_c), .CO(n17273));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_8_lut (.I0(GND_net), .I1(n843_adj_567[5]), 
            .I2(n129_c), .I3(n17271), .O(n842_adj_573[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_8 (.CI(n17271), .I0(n843_adj_567[5]), 
            .I1(n129_c), .CO(n17272));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_7_lut (.I0(GND_net), .I1(n843_adj_567[4]), 
            .I2(n129_c), .I3(n17270), .O(n842_adj_573[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_7 (.CI(n17270), .I0(n843_adj_567[4]), 
            .I1(n129_c), .CO(n17271));
    SB_LUT4 i1_2_lut_adj_128 (.I0(\Product_mul_temp[26] ), .I1(Error_sub_temp[29]), 
            .I2(GND_net), .I3(GND_net), .O(n789_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_2_lut_adj_128.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_6_lut (.I0(GND_net), .I1(n843_adj_567[3]), 
            .I2(n129_c), .I3(n17269), .O(n842_adj_573[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_6 (.CI(n17269), .I0(n843_adj_567[3]), 
            .I1(n129_c), .CO(n17270));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_5_lut (.I0(GND_net), .I1(n843_adj_567[2]), 
            .I2(n129_c), .I3(n17268), .O(n842_adj_573[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_5 (.CI(n17268), .I0(n843_adj_567[2]), 
            .I1(n129_c), .CO(n17269));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_4_lut (.I0(GND_net), .I1(n843_adj_567[1]), 
            .I2(n129_c), .I3(n17267), .O(n842_adj_573[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_4 (.CI(n17267), .I0(n843_adj_567[1]), 
            .I1(n129_c), .CO(n17268));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_3_lut (.I0(GND_net), .I1(n843_adj_567[0]), 
            .I2(n129_c), .I3(n17266), .O(n842_adj_573[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_3 (.CI(n17266), .I0(n843_adj_567[0]), 
            .I1(n129_c), .CO(n17267));
    SB_LUT4 paramCurrentControlP_15__I_0_add_571_2_lut (.I0(GND_net), .I1(n132_c), 
            .I2(n129_c), .I3(GND_net), .O(n842_adj_573[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_571_2 (.CI(GND_net), .I0(n132_c), 
            .I1(n129_c), .CO(n17266));
    SB_LUT4 add_559_33_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[31]), 
            .I3(n16003), .O(Saturate_out1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_32_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[30]), 
            .I3(n16002), .O(\Add_add_temp[34] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_32 (.CI(n16002), .I0(Switch_out1[31]), .I1(currentControlITerm[30]), 
            .CO(n16003));
    SB_LUT4 add_559_31_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[29]), 
            .I3(n16001), .O(\Add_add_temp[33] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_31 (.CI(n16001), .I0(Switch_out1[31]), .I1(currentControlITerm[29]), 
            .CO(n16002));
    SB_LUT4 add_559_30_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[28]), 
            .I3(n16000), .O(\Add_add_temp[32] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_30 (.CI(n16000), .I0(Switch_out1[31]), .I1(currentControlITerm[28]), 
            .CO(n16001));
    SB_LUT4 add_559_29_lut (.I0(GND_net), .I1(Switch_out1[31]), .I2(currentControlITerm[27]), 
            .I3(n15999), .O(\Add_add_temp[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_29 (.CI(n15999), .I0(Switch_out1[31]), .I1(currentControlITerm[27]), 
            .CO(n16000));
    SB_LUT4 add_559_28_lut (.I0(GND_net), .I1(Switch_out1[30]), .I2(currentControlITerm[26]), 
            .I3(n15998), .O(\Add_add_temp[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_28 (.CI(n15998), .I0(Switch_out1[30]), .I1(currentControlITerm[26]), 
            .CO(n15999));
    SB_LUT4 add_559_27_lut (.I0(GND_net), .I1(Switch_out1[29]), .I2(currentControlITerm[25]), 
            .I3(n15997), .O(\Add_add_temp[29] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_27 (.CI(n15997), .I0(Switch_out1[29]), .I1(currentControlITerm[25]), 
            .CO(n15998));
    SB_LUT4 add_559_26_lut (.I0(GND_net), .I1(Switch_out1[28]), .I2(currentControlITerm[24]), 
            .I3(n15996), .O(\Add_add_temp[28] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_26 (.CI(n15996), .I0(Switch_out1[28]), .I1(currentControlITerm[24]), 
            .CO(n15997));
    SB_LUT4 add_559_25_lut (.I0(GND_net), .I1(Switch_out1[27]), .I2(currentControlITerm[23]), 
            .I3(n15995), .O(\Add_add_temp[27] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_25 (.CI(n15995), .I0(Switch_out1[27]), .I1(currentControlITerm[23]), 
            .CO(n15996));
    SB_LUT4 add_559_24_lut (.I0(GND_net), .I1(Switch_out1[26]), .I2(currentControlITerm[22]), 
            .I3(n15994), .O(\Add_add_temp[26] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_24 (.CI(n15994), .I0(Switch_out1[26]), .I1(currentControlITerm[22]), 
            .CO(n15995));
    SB_LUT4 add_559_23_lut (.I0(GND_net), .I1(Switch_out1[25]), .I2(currentControlITerm[21]), 
            .I3(n15993), .O(\Add_add_temp[25] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_23 (.CI(n15993), .I0(Switch_out1[25]), .I1(currentControlITerm[21]), 
            .CO(n15994));
    SB_LUT4 add_559_22_lut (.I0(GND_net), .I1(Switch_out1[24]), .I2(currentControlITerm[20]), 
            .I3(n15992), .O(\Add_add_temp[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_22 (.CI(n15992), .I0(Switch_out1[24]), .I1(currentControlITerm[20]), 
            .CO(n15993));
    SB_LUT4 add_559_21_lut (.I0(GND_net), .I1(Switch_out1[23]), .I2(currentControlITerm[19]), 
            .I3(n15991), .O(\Add_add_temp[23] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_21 (.CI(n15991), .I0(Switch_out1[23]), .I1(currentControlITerm[19]), 
            .CO(n15992));
    SB_LUT4 add_559_20_lut (.I0(GND_net), .I1(Switch_out1[22]), .I2(currentControlITerm[18]), 
            .I3(n15990), .O(\Add_add_temp[22] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_20 (.CI(n15990), .I0(Switch_out1[22]), .I1(currentControlITerm[18]), 
            .CO(n15991));
    SB_LUT4 add_559_19_lut (.I0(GND_net), .I1(Switch_out1[21]), .I2(currentControlITerm[17]), 
            .I3(n15989), .O(\Add_add_temp[21] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_19 (.CI(n15989), .I0(Switch_out1[21]), .I1(currentControlITerm[17]), 
            .CO(n15990));
    SB_LUT4 add_559_18_lut (.I0(GND_net), .I1(Switch_out1[20]), .I2(currentControlITerm[16]), 
            .I3(n15988), .O(\Add_add_temp[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_18 (.CI(n15988), .I0(Switch_out1[20]), .I1(currentControlITerm[16]), 
            .CO(n15989));
    SB_LUT4 add_559_17_lut (.I0(GND_net), .I1(Switch_out1[19]), .I2(currentControlITerm[15]), 
            .I3(n15987), .O(\Add_add_temp[19] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_17 (.CI(n15987), .I0(Switch_out1[19]), .I1(currentControlITerm[15]), 
            .CO(n15988));
    SB_LUT4 add_559_16_lut (.I0(GND_net), .I1(Switch_out1[18]), .I2(currentControlITerm[14]), 
            .I3(n15986), .O(\Add_add_temp[18] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_16 (.CI(n15986), .I0(Switch_out1[18]), .I1(currentControlITerm[14]), 
            .CO(n15987));
    SB_LUT4 add_559_15_lut (.I0(GND_net), .I1(Switch_out1[17]), .I2(currentControlITerm[13]), 
            .I3(n15985), .O(\Add_add_temp[17] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_15 (.CI(n15985), .I0(Switch_out1[17]), .I1(currentControlITerm[13]), 
            .CO(n15986));
    SB_LUT4 add_559_14_lut (.I0(GND_net), .I1(Switch_out1[16]), .I2(currentControlITerm[12]), 
            .I3(n15984), .O(\Add_add_temp[16] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_14 (.CI(n15984), .I0(Switch_out1[16]), .I1(currentControlITerm[12]), 
            .CO(n15985));
    SB_LUT4 add_559_13_lut (.I0(GND_net), .I1(Switch_out1[15]), .I2(currentControlITerm[11]), 
            .I3(n15983), .O(\Add_add_temp[15] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_13 (.CI(n15983), .I0(Switch_out1[15]), .I1(currentControlITerm[11]), 
            .CO(n15984));
    SB_LUT4 add_559_12_lut (.I0(GND_net), .I1(Switch_out1[14]), .I2(currentControlITerm[10]), 
            .I3(n15982), .O(\Add_add_temp[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_12 (.CI(n15982), .I0(Switch_out1[14]), .I1(currentControlITerm[10]), 
            .CO(n15983));
    SB_LUT4 add_559_11_lut (.I0(GND_net), .I1(Switch_out1[13]), .I2(currentControlITerm[9]), 
            .I3(n15981), .O(\Add_add_temp[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_11 (.CI(n15981), .I0(Switch_out1[13]), .I1(currentControlITerm[9]), 
            .CO(n15982));
    SB_LUT4 add_559_10_lut (.I0(GND_net), .I1(Switch_out1[12]), .I2(currentControlITerm[8]), 
            .I3(n15980), .O(\Add_add_temp[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_10 (.CI(n15980), .I0(Switch_out1[12]), .I1(currentControlITerm[8]), 
            .CO(n15981));
    SB_LUT4 add_559_9_lut (.I0(GND_net), .I1(Switch_out1[11]), .I2(preSatVoltage[0]), 
            .I3(n15979), .O(\Add_add_temp[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_9 (.CI(n15979), .I0(Switch_out1[11]), .I1(preSatVoltage[0]), 
            .CO(n15980));
    SB_LUT4 add_559_8_lut (.I0(GND_net), .I1(Switch_out1[10]), .I2(currentControlITerm[6]), 
            .I3(n15978), .O(\Add_add_temp[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_8 (.CI(n15978), .I0(Switch_out1[10]), .I1(currentControlITerm[6]), 
            .CO(n15979));
    SB_LUT4 add_559_7_lut (.I0(GND_net), .I1(Switch_out1[9]), .I2(currentControlITerm[5]), 
            .I3(n15977), .O(\Add_add_temp[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_7 (.CI(n15977), .I0(Switch_out1[9]), .I1(currentControlITerm[5]), 
            .CO(n15978));
    SB_LUT4 add_559_6_lut (.I0(GND_net), .I1(Switch_out1[8]), .I2(currentControlITerm[4]), 
            .I3(n15976), .O(\Add_add_temp[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_6 (.CI(n15976), .I0(Switch_out1[8]), .I1(currentControlITerm[4]), 
            .CO(n15977));
    SB_LUT4 add_559_5_lut (.I0(GND_net), .I1(Switch_out1[7]), .I2(currentControlITerm[3]), 
            .I3(n15975), .O(\Add_add_temp[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_5 (.CI(n15975), .I0(Switch_out1[7]), .I1(currentControlITerm[3]), 
            .CO(n15976));
    SB_LUT4 add_559_4_lut (.I0(GND_net), .I1(Switch_out1[6]), .I2(currentControlITerm[2]), 
            .I3(n15974), .O(\Add_add_temp[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_9 (.CI(n17772), .I0(n836_adj_565[6]), 
            .I1(n123_c), .CO(n17773));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_8_lut (.I0(GND_net), .I1(n836_adj_565[5]), 
            .I2(n120_c), .I3(n17771), .O(n835_adj_564[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_8 (.CI(n17771), .I0(n836_adj_565[5]), 
            .I1(n120_c), .CO(n17772));
    SB_LUT4 i1_4_lut_adj_129 (.I0(n789_c), .I1(n142), .I2(n19269), .I3(n19273), 
            .O(n791));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_adj_129.LUT_INIT = 16'heca8;
    SB_CARRY Error_sub_temp_31__I_0_add_562_6 (.CI(n17739), .I0(n834_adj_574[3]), 
            .I1(n114_c), .CO(n17740));
    SB_CARRY add_4257_6 (.CI(n17715), .I0(n836_adj_565[14]), .I1(n751), 
            .CO(n17716));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_5_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[2]), .I2(n111_c), .I3(n17738), .O(Switch_out1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Error_sub_temp_31__I_0_add_564_7_lut (.I0(GND_net), .I1(n836_adj_565[4]), 
            .I2(n117_c), .I3(n17770), .O(n835_adj_564[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_7 (.CI(n17770), .I0(n836_adj_565[4]), 
            .I1(n117_c), .CO(n17771));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_12_lut (.I0(GND_net), .I1(n838_adj_571[9]), 
            .I2(n132_c), .I3(n17805), .O(n837_adj_572[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_16 (.CI(n17824), .I0(n839_adj_570[13]), 
            .I1(n146), .CO(n763));
    SB_LUT4 add_4257_5_lut (.I0(Not_Equal_relop1_N_201), .I1(n835_adj_564[14]), 
            .I2(n747), .I3(n17714), .O(Switch_out1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_15_lut (.I0(GND_net), .I1(n839_adj_570[12]), 
            .I2(n141), .I3(n17823), .O(n838_adj_571[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_11 (.CI(n17649), .I0(n841[8]), 
            .I1(n123_c), .CO(n17650));
    SB_CARRY add_4257_5 (.CI(n17714), .I0(n835_adj_564[14]), .I1(n747), 
            .CO(n17715));
    SB_CARRY Error_sub_temp_31__I_0_add_562_5 (.CI(n17738), .I0(n834_adj_574[2]), 
            .I1(n111_c), .CO(n17739));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_4_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[1]), .I2(n108_c), .I3(n17737), .O(Switch_out1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4257_4_lut (.I0(Not_Equal_relop1_N_201), .I1(n834_adj_574[14]), 
            .I2(n743), .I3(n17713), .O(Switch_out1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4257_4 (.CI(n17713), .I0(n834_adj_574[14]), .I1(n743), 
            .CO(n17714));
    SB_CARRY add_3099_12 (.CI(n17515), .I0(n842_adj_573[14]), .I1(n775_adj_357), 
            .CO(n17516));
    SB_CARRY Error_sub_temp_31__I_0_add_567_15 (.CI(n17823), .I0(n839_adj_570[12]), 
            .I1(n141), .CO(n17824));
    SB_CARRY Error_sub_temp_31__I_0_add_566_12 (.CI(n17805), .I0(n838_adj_571[9]), 
            .I1(n132_c), .CO(n17806));
    SB_CARRY add_559_4 (.CI(n15974), .I0(Switch_out1[6]), .I1(currentControlITerm[2]), 
            .CO(n15975));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_6_lut (.I0(GND_net), .I1(n836_adj_565[3]), 
            .I2(n114_c), .I3(n17769), .O(n835_adj_564[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4257_3_lut (.I0(Not_Equal_relop1_N_201), .I1(n833_adj_575[14]), 
            .I2(n8265), .I3(n17712), .O(Switch_out1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_564_6 (.CI(n17769), .I0(n836_adj_565[3]), 
            .I1(n114_c), .CO(n17770));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_11_lut (.I0(GND_net), .I1(n838_adj_571[8]), 
            .I2(n129_c), .I3(n17804), .O(n837_adj_572[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_14_lut (.I0(GND_net), .I1(n839_adj_570[11]), 
            .I2(n138_c), .I3(n17822), .O(n838_adj_571[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_4 (.CI(n17737), .I0(n834_adj_574[1]), 
            .I1(n108_c), .CO(n17738));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_5_lut (.I0(GND_net), .I1(n836_adj_565[2]), 
            .I2(n111_c), .I3(n17768), .O(n835_adj_564[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_11_lut (.I0(GND_net), .I1(n841[14]), .I2(n771), .I3(n17514), 
            .O(Proportional_Gain_mul_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_5 (.CI(n17768), .I0(n836_adj_565[2]), 
            .I1(n111_c), .CO(n17769));
    SB_CARRY Error_sub_temp_31__I_0_add_566_11 (.CI(n17804), .I0(n838_adj_571[8]), 
            .I1(n129_c), .CO(n17805));
    SB_LUT4 add_559_3_lut (.I0(GND_net), .I1(Switch_out1[5]), .I2(currentControlITerm[1]), 
            .I3(n15973), .O(\Add_add_temp[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_14 (.CI(n17822), .I0(n839_adj_570[11]), 
            .I1(n138_c), .CO(n17823));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_5_lut (.I0(GND_net), .I1(n835_adj_564[2]), 
            .I2(n111_c), .I3(n17753), .O(n834_adj_574[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_566_10_lut (.I0(GND_net), .I1(n838_adj_571[7]), 
            .I2(n126_c), .I3(n17803), .O(n837_adj_572[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_10 (.CI(n17803), .I0(n838_adj_571[7]), 
            .I1(n126_c), .CO(n17804));
    SB_LUT4 paramCurrentControlP_15__I_0_i542_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(\Error_sub_temp[31] ), .I2(GND_net), .I3(GND_net), .O(n796));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i542_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_9 (.CI(n17557), .I0(n835[6]), 
            .I1(n105_c), .CO(n17558));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_14_lut (.I0(GND_net), .I1(n835[11]), 
            .I2(n105_c), .I3(n17562), .O(n834[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_11 (.CI(n17514), .I0(n841[14]), .I1(n771), .CO(n17515));
    SB_CARRY paramCurrentControlP_15__I_0_add_563_14 (.CI(n17562), .I0(n835[11]), 
            .I1(n105_c), .CO(n17563));
    SB_LUT4 i6572_2_lut (.I0(n833_adj_575[13]), .I1(\Error_sub_temp[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n8265));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(92[30:64])
    defparam i6572_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Error_sub_temp_31__I_0_add_572_4 (.CI(n17898), .I0(n844[1]), 
            .I1(n108_c), .CO(n17899));
    SB_LUT4 paramCurrentControlP_15__I_0_i37_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[17]), .I2(GND_net), .I3(GND_net), .O(n102_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i37_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_13_lut (.I0(GND_net), .I1(n839_adj_570[10]), 
            .I2(n135_c), .I3(n17821), .O(n838_adj_571[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_3 (.CI(n15973), .I0(Switch_out1[5]), .I1(currentControlITerm[1]), 
            .CO(n15974));
    SB_LUT4 add_559_2_lut (.I0(GND_net), .I1(Switch_out1[4]), .I2(currentControlITerm[0]), 
            .I3(GND_net), .O(\Add_add_temp[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_572_6_lut (.I0(GND_net), .I1(n844[3]), 
            .I2(n114_c), .I3(n17900), .O(n843[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_566_9_lut (.I0(GND_net), .I1(n838_adj_571[6]), 
            .I2(n123_c), .I3(n17802), .O(n837_adj_572[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_564_4_lut (.I0(GND_net), .I1(n836_adj_565[1]), 
            .I2(n108_c), .I3(n17767), .O(n835_adj_564[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_9 (.CI(n17802), .I0(n838_adj_571[6]), 
            .I1(n123_c), .CO(n17803));
    SB_CARRY Error_sub_temp_31__I_0_add_564_4 (.CI(n17767), .I0(n836_adj_565[1]), 
            .I1(n108_c), .CO(n17768));
    SB_LUT4 add_3099_10_lut (.I0(GND_net), .I1(n840[14]), .I2(n767_adj_382), 
            .I3(n17513), .O(Proportional_Gain_mul_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_10 (.CI(n17513), .I0(n840[14]), .I1(n767_adj_382), 
            .CO(n17514));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_3_lut (.I0(GND_net), .I1(n836_adj_565[0]), 
            .I2(n105_c), .I3(n17766), .O(n835_adj_564[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_9_lut (.I0(GND_net), .I1(n839[14]), .I2(n763_adj_386), 
            .I3(n17512), .O(Proportional_Gain_mul_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_6 (.CI(n17900), .I0(n844[3]), 
            .I1(n114_c), .CO(n17901));
    SB_CARRY Error_sub_temp_31__I_0_add_564_3 (.CI(n17766), .I0(n836_adj_565[0]), 
            .I1(n105_c), .CO(n17767));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_5_lut (.I0(GND_net), .I1(n844[2]), 
            .I2(n111_c), .I3(n17899), .O(n843[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_9 (.CI(n17512), .I0(n839[14]), .I1(n763_adj_386), 
            .CO(n17513));
    SB_CARRY add_559_2 (.CI(GND_net), .I0(Switch_out1[4]), .I1(currentControlITerm[0]), 
            .CO(n15973));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_3_lut (.I0(GND_net), .I1(n844[0]), 
            .I2(n105_c), .I3(n17897), .O(n843[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_10 (.CI(n17573), .I0(n836[7]), 
            .I1(n108_c), .CO(n17574));
    SB_CARRY Error_sub_temp_31__I_0_add_572_3 (.CI(n17897), .I0(n844[0]), 
            .I1(n105_c), .CO(n17898));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n843[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_9_lut (.I0(GND_net), .I1(n836[6]), 
            .I2(n108_c), .I3(n17572), .O(n835[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17897));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_16_lut (.I0(GND_net), .I1(n843[13]), 
            .I2(n146), .I3(n17895), .O(n842[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_16 (.CI(n17895), .I0(n843[13]), 
            .I1(n146), .CO(n779));
    SB_CARRY paramCurrentControlP_15__I_0_add_564_9 (.CI(n17572), .I0(n836[6]), 
            .I1(n108_c), .CO(n17573));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_8_lut (.I0(GND_net), .I1(n836[5]), 
            .I2(n108_c), .I3(n17571), .O(n835[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_8 (.CI(n17571), .I0(n836[5]), 
            .I1(n108_c), .CO(n17572));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_7_lut (.I0(GND_net), .I1(n836[4]), 
            .I2(n108_c), .I3(n17570), .O(n835[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_13 (.CI(n17821), .I0(n839_adj_570[10]), 
            .I1(n135_c), .CO(n17822));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_15_lut (.I0(GND_net), .I1(n843[12]), 
            .I2(n141), .I3(n17894), .O(n842[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF currentControlITerm_i9 (.Q(currentControlITerm[9]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14328));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 paramCurrentControlP_15__I_0_i59_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[28]), .I2(GND_net), .I3(GND_net), .O(n135_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_7 (.CI(n17570), .I0(n836[4]), 
            .I1(n108_c), .CO(n17571));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_6_lut (.I0(GND_net), .I1(n836[3]), 
            .I2(n108_c), .I3(n17569), .O(n835[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF currentControlITerm_i8 (.Q(currentControlITerm[8]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14327));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i7 (.Q(preSatVoltage[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14326));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_CARRY paramCurrentControlP_15__I_0_add_564_6 (.CI(n17569), .I0(n836[3]), 
            .I1(n108_c), .CO(n17570));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_5_lut (.I0(GND_net), .I1(n836[2]), 
            .I2(n108_c), .I3(n17568), .O(n835[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF currentControlITerm_i3 (.Q(currentControlITerm[3]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14322));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_CARRY paramCurrentControlP_15__I_0_add_562_15 (.CI(n17548), .I0(n834[12]), 
            .I1(n102_c), .CO(n17549));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_8_lut (.I0(GND_net), .I1(n835[5]), 
            .I2(n105_c), .I3(n17556), .O(n834[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_7 (.CI(n17585), .I0(n837[4]), 
            .I1(n111_c), .CO(n17586));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_8_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n785_c), .I3(n18172), .O(n844_adj_566[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_8 (.CI(n18172), .I0(n845[3]), 
            .I1(n785_c), .CO(n787));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_7_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n135_c), .I3(n18171), .O(n844_adj_566[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_7 (.CI(n18171), .I0(n845[3]), 
            .I1(n135_c), .CO(n18172));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_6_lut (.I0(GND_net), .I1(n845[3]), 
            .I2(n135_c), .I3(n18170), .O(n844_adj_566[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_6 (.CI(n18170), .I0(n845[3]), 
            .I1(n135_c), .CO(n18171));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_5_lut (.I0(GND_net), .I1(n845[2]), 
            .I2(n135_c), .I3(n18169), .O(n844_adj_566[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_5 (.CI(n18169), .I0(n845[2]), 
            .I1(n135_c), .CO(n18170));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_4_lut (.I0(GND_net), .I1(n845[1]), 
            .I2(n135_c), .I3(n18168), .O(n844_adj_566[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_4 (.CI(n18168), .I0(n845[1]), 
            .I1(n135_c), .CO(n18169));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_3_lut (.I0(GND_net), .I1(n845[0]), 
            .I2(n135_c), .I3(n18167), .O(n844_adj_566[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_3 (.CI(n18167), .I0(n845[0]), 
            .I1(n135_c), .CO(n18168));
    SB_LUT4 paramCurrentControlP_15__I_0_add_573_2_lut (.I0(GND_net), .I1(n138_c), 
            .I2(n135_c), .I3(GND_net), .O(n844_adj_566[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_573_2 (.CI(GND_net), .I0(n138_c), 
            .I1(n135_c), .CO(n18167));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_8_lut (.I0(GND_net), .I1(n838_adj_571[5]), 
            .I2(n120_c), .I3(n17801), .O(n837_adj_572[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_8_lut (.I0(GND_net), .I1(n838[14]), .I2(n759), .I3(n17511), 
            .O(Proportional_Gain_mul_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_8 (.CI(n17511), .I0(n838[14]), .I1(n759), .CO(n17512));
    SB_LUT4 add_3099_7_lut (.I0(GND_net), .I1(n837[14]), .I2(n755_adj_404), 
            .I3(n17510), .O(Proportional_Gain_mul_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_7 (.CI(n17510), .I0(n837[14]), .I1(n755_adj_404), 
            .CO(n17511));
    SB_LUT4 add_3099_6_lut (.I0(GND_net), .I1(n836[14]), .I2(n751_adj_406), 
            .I3(n17509), .O(Proportional_Gain_mul_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_6 (.CI(n17509), .I0(n836[14]), .I1(n751_adj_406), 
            .CO(n17510));
    SB_LUT4 add_3099_5_lut (.I0(GND_net), .I1(n835[14]), .I2(n747_adj_408), 
            .I3(n17508), .O(Proportional_Gain_mul_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_5 (.CI(n17508), .I0(n835[14]), .I1(n747_adj_408), 
            .CO(n17509));
    SB_LUT4 add_3099_4_lut (.I0(GND_net), .I1(n834[14]), .I2(n743_adj_410), 
            .I3(n17507), .O(Proportional_Gain_mul_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_4 (.CI(n17507), .I0(n834[14]), .I1(n743_adj_410), 
            .CO(n17508));
    SB_LUT4 add_3099_3_lut (.I0(GND_net), .I1(n833[14]), .I2(n739), .I3(n17506), 
            .O(Proportional_Gain_mul_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_3 (.CI(n17506), .I0(n833[14]), .I1(n739), .CO(n17507));
    SB_LUT4 add_3099_2_lut (.I0(GND_net), .I1(\Product_mul_temp[26] ), .I2(\Error_sub_temp[31] ), 
            .I3(n17505), .O(Proportional_Gain_mul_temp[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_2 (.CI(n17505), .I0(\Product_mul_temp[26] ), .I1(\Error_sub_temp[31] ), 
            .CO(n17506));
    SB_CARRY add_3099_1 (.CI(GND_net), .I0(n832[14]), .I1(n832[14]), .CO(n17505));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_12_lut (.I0(GND_net), .I1(n839_adj_570[9]), 
            .I2(n132_c), .I3(n17820), .O(n838_adj_571[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_15 (.CI(n17894), .I0(n843[12]), 
            .I1(n141), .CO(n17895));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_3_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[0]), .I2(n105_c), .I3(n17736), .O(Switch_out1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_10_lut (.I0(GND_net), .I1(n844_adj_566[5]), 
            .I2(n781_c), .I3(n18142), .O(n843_adj_567[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_10 (.CI(n18142), .I0(n844_adj_566[5]), 
            .I1(n781_c), .CO(n783_adj_349));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_9_lut (.I0(GND_net), .I1(n844_adj_566[5]), 
            .I2(n132_c), .I3(n18141), .O(n843_adj_567[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_9 (.CI(n18141), .I0(n844_adj_566[5]), 
            .I1(n132_c), .CO(n18142));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_8_lut (.I0(GND_net), .I1(n844_adj_566[5]), 
            .I2(n132_c), .I3(n18140), .O(n843_adj_567[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_8 (.CI(n18140), .I0(n844_adj_566[5]), 
            .I1(n132_c), .CO(n18141));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_7_lut (.I0(GND_net), .I1(n844_adj_566[4]), 
            .I2(n132_c), .I3(n18139), .O(n843_adj_567[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_7 (.CI(n18139), .I0(n844_adj_566[4]), 
            .I1(n132_c), .CO(n18140));
    SB_CARRY Error_sub_temp_31__I_0_add_567_12 (.CI(n17820), .I0(n839_adj_570[9]), 
            .I1(n132_c), .CO(n17821));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_6_lut (.I0(GND_net), .I1(n844_adj_566[3]), 
            .I2(n132_c), .I3(n18138), .O(n843_adj_567[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_6 (.CI(n18138), .I0(n844_adj_566[3]), 
            .I1(n132_c), .CO(n18139));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_5_lut (.I0(GND_net), .I1(n844_adj_566[2]), 
            .I2(n132_c), .I3(n18137), .O(n843_adj_567[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_5 (.CI(n18137), .I0(n844_adj_566[2]), 
            .I1(n132_c), .CO(n18138));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_4_lut (.I0(GND_net), .I1(n844_adj_566[1]), 
            .I2(n132_c), .I3(n18136), .O(n843_adj_567[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_4 (.CI(n18136), .I0(n844_adj_566[1]), 
            .I1(n132_c), .CO(n18137));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_3_lut (.I0(GND_net), .I1(n844_adj_566[0]), 
            .I2(n132_c), .I3(n18135), .O(n843_adj_567[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_3 (.CI(n18135), .I0(n844_adj_566[0]), 
            .I1(n132_c), .CO(n18136));
    SB_LUT4 paramCurrentControlP_15__I_0_add_572_2_lut (.I0(GND_net), .I1(n135_c), 
            .I2(n132_c), .I3(GND_net), .O(n843_adj_567[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_572_2 (.CI(GND_net), .I0(n135_c), 
            .I1(n132_c), .CO(n18135));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_14_lut (.I0(GND_net), .I1(n842_adj_573[9]), 
            .I2(n773_c), .I3(n18133), .O(n841[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_14 (.CI(n18133), .I0(n842_adj_573[9]), 
            .I1(n773_c), .CO(n775_adj_357));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_13_lut (.I0(GND_net), .I1(n842_adj_573[9]), 
            .I2(n126_c), .I3(n18132), .O(n841[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_13 (.CI(n18132), .I0(n842_adj_573[9]), 
            .I1(n126_c), .CO(n18133));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_12_lut (.I0(GND_net), .I1(n842_adj_573[9]), 
            .I2(n126_c), .I3(n18131), .O(n841[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_12 (.CI(n18131), .I0(n842_adj_573[9]), 
            .I1(n126_c), .CO(n18132));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_11_lut (.I0(GND_net), .I1(n842_adj_573[8]), 
            .I2(n126_c), .I3(n18130), .O(n841[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_11 (.CI(n18130), .I0(n842_adj_573[8]), 
            .I1(n126_c), .CO(n18131));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_10_lut (.I0(GND_net), .I1(n842_adj_573[7]), 
            .I2(n126_c), .I3(n18129), .O(n841[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_10 (.CI(n18129), .I0(n842_adj_573[7]), 
            .I1(n126_c), .CO(n18130));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_9_lut (.I0(GND_net), .I1(n842_adj_573[6]), 
            .I2(n126_c), .I3(n18128), .O(n841[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_9 (.CI(n18128), .I0(n842_adj_573[6]), 
            .I1(n126_c), .CO(n18129));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_8_lut (.I0(GND_net), .I1(n842_adj_573[5]), 
            .I2(n126_c), .I3(n18127), .O(n841[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_8 (.CI(n18127), .I0(n842_adj_573[5]), 
            .I1(n126_c), .CO(n18128));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_7_lut (.I0(GND_net), .I1(n842_adj_573[4]), 
            .I2(n126_c), .I3(n18126), .O(n841[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_7 (.CI(n18126), .I0(n842_adj_573[4]), 
            .I1(n126_c), .CO(n18127));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_6_lut (.I0(GND_net), .I1(n842_adj_573[3]), 
            .I2(n126_c), .I3(n18125), .O(n841[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_6 (.CI(n18125), .I0(n842_adj_573[3]), 
            .I1(n126_c), .CO(n18126));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_5_lut (.I0(GND_net), .I1(n842_adj_573[2]), 
            .I2(n126_c), .I3(n18124), .O(n841[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_5 (.CI(n18124), .I0(n842_adj_573[2]), 
            .I1(n126_c), .CO(n18125));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_4_lut (.I0(GND_net), .I1(n842_adj_573[1]), 
            .I2(n126_c), .I3(n18123), .O(n841[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_4 (.CI(n18123), .I0(n842_adj_573[1]), 
            .I1(n126_c), .CO(n18124));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_3_lut (.I0(GND_net), .I1(n842_adj_573[0]), 
            .I2(n126_c), .I3(n18122), .O(n841[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_3 (.CI(n18122), .I0(n842_adj_573[0]), 
            .I1(n126_c), .CO(n18123));
    SB_LUT4 paramCurrentControlP_15__I_0_add_570_2_lut (.I0(GND_net), .I1(n129_c), 
            .I2(n126_c), .I3(GND_net), .O(n841[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_570_2 (.CI(GND_net), .I0(n129_c), 
            .I1(n126_c), .CO(n18122));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_16_lut (.I0(GND_net), .I1(n793), 
            .I2(n146), .I3(n17955), .O(n846[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_16 (.CI(n17955), .I0(n793), 
            .I1(n146), .CO(n795));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_15_lut (.I0(GND_net), .I1(n789_c), 
            .I2(n141), .I3(n17954), .O(n846[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_15 (.CI(n17954), .I0(n789_c), 
            .I1(n141), .CO(n17955));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_14_lut (.I0(GND_net), .I1(n785_c), 
            .I2(n138_c), .I3(n17953), .O(n846[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_14 (.CI(n17953), .I0(n785_c), 
            .I1(n138_c), .CO(n17954));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_13_lut (.I0(GND_net), .I1(n781_c), 
            .I2(n135_c), .I3(n17952), .O(n846[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_13 (.CI(n17952), .I0(n781_c), 
            .I1(n135_c), .CO(n17953));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_12_lut (.I0(GND_net), .I1(n777_c), 
            .I2(n132_c), .I3(n17951), .O(n846[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_12 (.CI(n17951), .I0(n777_c), 
            .I1(n132_c), .CO(n17952));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_11_lut (.I0(GND_net), .I1(n773_c), 
            .I2(n129_c), .I3(n17950), .O(n846[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_11 (.CI(n17950), .I0(n773_c), 
            .I1(n129_c), .CO(n17951));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_10_lut (.I0(GND_net), .I1(n769_c), 
            .I2(n126_c), .I3(n17949), .O(n846[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_10 (.CI(n17949), .I0(n769_c), 
            .I1(n126_c), .CO(n17950));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_9_lut (.I0(GND_net), .I1(n765_c), 
            .I2(n123_c), .I3(n17948), .O(n846[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_9 (.CI(n17948), .I0(n765_c), 
            .I1(n123_c), .CO(n17949));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_8_lut (.I0(GND_net), .I1(n761_c), 
            .I2(n120_c), .I3(n17947), .O(n846[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_8 (.CI(n17947), .I0(n761_c), 
            .I1(n120_c), .CO(n17948));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_7_lut (.I0(GND_net), .I1(n757_c), 
            .I2(n117_c), .I3(n17946), .O(n846[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_7 (.CI(n17946), .I0(n757_c), 
            .I1(n117_c), .CO(n17947));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_6_lut (.I0(GND_net), .I1(n753_c), 
            .I2(n114_c), .I3(n17945), .O(n846[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_6 (.CI(n17945), .I0(n753_c), 
            .I1(n114_c), .CO(n17946));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_5_lut (.I0(GND_net), .I1(n749_c), 
            .I2(n111_c), .I3(n17944), .O(n846[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_5 (.CI(n17944), .I0(n749_c), 
            .I1(n111_c), .CO(n17945));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_4_lut (.I0(GND_net), .I1(n745_c), 
            .I2(n108_c), .I3(n17943), .O(n846[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_4 (.CI(n17943), .I0(n745_c), 
            .I1(n108_c), .CO(n17944));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_3_lut (.I0(GND_net), .I1(n741_c), 
            .I2(n105_c), .I3(n17942), .O(n846[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_3 (.CI(n17942), .I0(n741_c), 
            .I1(n105_c), .CO(n17943));
    SB_LUT4 Error_sub_temp_31__I_0_add_575_2_lut (.I0(GND_net), .I1(n737_c), 
            .I2(n102_c), .I3(GND_net), .O(n846[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_575_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_575_2 (.CI(GND_net), .I0(n737_c), 
            .I1(n102_c), .CO(n17942));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_16_lut (.I0(GND_net), .I1(n846[13]), 
            .I2(n146), .I3(n17940), .O(n845_adj_576[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_16 (.CI(n17940), .I0(n846[13]), 
            .I1(n146), .CO(n791_adj_416));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_15_lut (.I0(GND_net), .I1(n846[12]), 
            .I2(n141), .I3(n17939), .O(n845_adj_576[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_15 (.CI(n17939), .I0(n846[12]), 
            .I1(n141), .CO(n17940));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_14_lut (.I0(GND_net), .I1(n846[11]), 
            .I2(n138_c), .I3(n17938), .O(n845_adj_576[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_14 (.CI(n17938), .I0(n846[11]), 
            .I1(n138_c), .CO(n17939));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_13_lut (.I0(GND_net), .I1(n846[10]), 
            .I2(n135_c), .I3(n17937), .O(n845_adj_576[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_13 (.CI(n17937), .I0(n846[10]), 
            .I1(n135_c), .CO(n17938));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_12_lut (.I0(GND_net), .I1(n846[9]), 
            .I2(n132_c), .I3(n17936), .O(n845_adj_576[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_12 (.CI(n17936), .I0(n846[9]), 
            .I1(n132_c), .CO(n17937));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_11_lut (.I0(GND_net), .I1(n846[8]), 
            .I2(n129_c), .I3(n17935), .O(n845_adj_576[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_11 (.CI(n17935), .I0(n846[8]), 
            .I1(n129_c), .CO(n17936));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_10_lut (.I0(GND_net), .I1(n846[7]), 
            .I2(n126_c), .I3(n17934), .O(n845_adj_576[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_10 (.CI(n17934), .I0(n846[7]), 
            .I1(n126_c), .CO(n17935));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_9_lut (.I0(GND_net), .I1(n846[6]), 
            .I2(n123_c), .I3(n17933), .O(n845_adj_576[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_9 (.CI(n17933), .I0(n846[6]), 
            .I1(n123_c), .CO(n17934));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_8_lut (.I0(GND_net), .I1(n846[5]), 
            .I2(n120_c), .I3(n17932), .O(n845_adj_576[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_8 (.CI(n17932), .I0(n846[5]), 
            .I1(n120_c), .CO(n17933));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_7_lut (.I0(GND_net), .I1(n846[4]), 
            .I2(n117_c), .I3(n17931), .O(n845_adj_576[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_7 (.CI(n17931), .I0(n846[4]), 
            .I1(n117_c), .CO(n17932));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_6_lut (.I0(GND_net), .I1(n846[3]), 
            .I2(n114_c), .I3(n17930), .O(n845_adj_576[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_6 (.CI(n17930), .I0(n846[3]), 
            .I1(n114_c), .CO(n17931));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_5_lut (.I0(GND_net), .I1(n846[2]), 
            .I2(n111_c), .I3(n17929), .O(n845_adj_576[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_5 (.CI(n17929), .I0(n846[2]), 
            .I1(n111_c), .CO(n17930));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_4_lut (.I0(GND_net), .I1(n846[1]), 
            .I2(n108_c), .I3(n17928), .O(n845_adj_576[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_4 (.CI(n17928), .I0(n846[1]), 
            .I1(n108_c), .CO(n17929));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_3_lut (.I0(GND_net), .I1(n846[0]), 
            .I2(n105_c), .I3(n17927), .O(n845_adj_576[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_3 (.CI(n17927), .I0(n846[0]), 
            .I1(n105_c), .CO(n17928));
    SB_LUT4 Error_sub_temp_31__I_0_add_574_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n845_adj_576[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_574_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_574_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17927));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_16_lut (.I0(GND_net), .I1(n845_adj_576[13]), 
            .I2(n146), .I3(n17925), .O(n844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_16 (.CI(n17925), .I0(n845_adj_576[13]), 
            .I1(n146), .CO(n787_adj_421));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_15_lut (.I0(GND_net), .I1(n845_adj_576[12]), 
            .I2(n141), .I3(n17924), .O(n844[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_15 (.CI(n17924), .I0(n845_adj_576[12]), 
            .I1(n141), .CO(n17925));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_14_lut (.I0(GND_net), .I1(n845_adj_576[11]), 
            .I2(n138_c), .I3(n17923), .O(n844[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_14 (.CI(n17923), .I0(n845_adj_576[11]), 
            .I1(n138_c), .CO(n17924));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_13_lut (.I0(GND_net), .I1(n845_adj_576[10]), 
            .I2(n135_c), .I3(n17922), .O(n844[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_13 (.CI(n17922), .I0(n845_adj_576[10]), 
            .I1(n135_c), .CO(n17923));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_10_lut (.I0(GND_net), .I1(n845_adj_576[7]), 
            .I2(n126_c), .I3(n17919), .O(n844[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_11 (.CI(n17920), .I0(n845_adj_576[8]), 
            .I1(n129_c), .CO(n17921));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_11_lut (.I0(GND_net), .I1(n845_adj_576[8]), 
            .I2(n129_c), .I3(n17920), .O(n844[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_8 (.CI(n17556), .I0(n835[5]), 
            .I1(n105_c), .CO(n17557));
    SB_CARRY Error_sub_temp_31__I_0_add_573_12 (.CI(n17921), .I0(n845_adj_576[9]), 
            .I1(n132_c), .CO(n17922));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_14_lut (.I0(GND_net), .I1(n843[11]), 
            .I2(n138_c), .I3(n17893), .O(n842[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_16_lut (.I0(GND_net), .I1(n836[13]), 
            .I2(n749_c), .I3(n17579), .O(n835[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_14 (.CI(n17893), .I0(n843[11]), 
            .I1(n138_c), .CO(n17894));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_13_lut (.I0(GND_net), .I1(n843[10]), 
            .I2(n135_c), .I3(n17892), .O(n842[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_5 (.CI(n17753), .I0(n835_adj_564[2]), 
            .I1(n111_c), .CO(n17754));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n835_adj_564[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_16 (.CI(n17579), .I0(n836[13]), 
            .I1(n749_c), .CO(n751_adj_406));
    SB_CARRY Error_sub_temp_31__I_0_add_566_8 (.CI(n17801), .I0(n838_adj_571[5]), 
            .I1(n120_c), .CO(n17802));
    SB_CARRY Error_sub_temp_31__I_0_add_571_13 (.CI(n17892), .I0(n843[10]), 
            .I1(n135_c), .CO(n17893));
    SB_CARRY Error_sub_temp_31__I_0_add_564_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17766));
    SB_CARRY add_4257_3 (.CI(n17712), .I0(n833_adj_575[14]), .I1(n8265), 
            .CO(n17713));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_7_lut (.I0(GND_net), .I1(n838_adj_571[4]), 
            .I2(n117_c), .I3(n17800), .O(n837_adj_572[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4257_2_lut (.I0(Not_Equal_relop1_N_201), .I1(\Error_sub_temp[31] ), 
            .I2(\Product_mul_temp[26] ), .I3(n17711), .O(Switch_out1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_11_lut (.I0(GND_net), .I1(n839_adj_570[8]), 
            .I2(n129_c), .I3(n17819), .O(n838_adj_571[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4257_2 (.CI(n17711), .I0(\Error_sub_temp[31] ), .I1(\Product_mul_temp[26] ), 
            .CO(n17712));
    SB_CARRY Error_sub_temp_31__I_0_add_567_11 (.CI(n17819), .I0(n839_adj_570[8]), 
            .I1(n129_c), .CO(n17820));
    SB_CARRY Error_sub_temp_31__I_0_add_566_7 (.CI(n17800), .I0(n838_adj_571[4]), 
            .I1(n117_c), .CO(n17801));
    SB_CARRY add_4257_1 (.CI(GND_net), .I0(n832_adj_577[14]), .I1(n832_adj_577[14]), 
            .CO(n17711));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_6_lut (.I0(GND_net), .I1(n838_adj_571[3]), 
            .I2(n114_c), .I3(n17799), .O(n837_adj_572[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_563_16_lut (.I0(GND_net), .I1(n835_adj_564[13]), 
            .I2(n146), .I3(n17764), .O(n834_adj_574[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_16 (.CI(n17764), .I0(n835_adj_564[13]), 
            .I1(n146), .CO(n747));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_10_lut (.I0(GND_net), .I1(n839_adj_570[7]), 
            .I2(n126_c), .I3(n17818), .O(n838_adj_571[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_10 (.CI(n17818), .I0(n839_adj_570[7]), 
            .I1(n126_c), .CO(n17819));
    SB_CARRY Error_sub_temp_31__I_0_add_562_3 (.CI(n17736), .I0(n834_adj_574[0]), 
            .I1(n105_c), .CO(n17737));
    SB_CARRY Error_sub_temp_31__I_0_add_562_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17736));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_9_lut (.I0(GND_net), .I1(n839_adj_570[6]), 
            .I2(n123_c), .I3(n17817), .O(n838_adj_571[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_5 (.CI(n17568), .I0(n836[2]), 
            .I1(n108_c), .CO(n17569));
    SB_CARRY Error_sub_temp_31__I_0_add_567_9 (.CI(n17817), .I0(n839_adj_570[6]), 
            .I1(n123_c), .CO(n17818));
    SB_CARRY Error_sub_temp_31__I_0_add_566_6 (.CI(n17799), .I0(n838_adj_571[3]), 
            .I1(n114_c), .CO(n17800));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_5_lut (.I0(GND_net), .I1(n838_adj_571[2]), 
            .I2(n111_c), .I3(n17798), .O(n837_adj_572[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_563_4_lut (.I0(GND_net), .I1(n835_adj_564[1]), 
            .I2(n108_c), .I3(n17752), .O(n834_adj_574[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_5 (.CI(n17798), .I0(n838_adj_571[2]), 
            .I1(n111_c), .CO(n17799));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_4_lut (.I0(GND_net), .I1(n838_adj_571[1]), 
            .I2(n108_c), .I3(n17797), .O(n837_adj_572[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_571_12_lut (.I0(GND_net), .I1(n843[9]), 
            .I2(n132_c), .I3(n17891), .O(n842[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_4 (.CI(n17752), .I0(n835_adj_564[1]), 
            .I1(n108_c), .CO(n17753));
    SB_CARRY Error_sub_temp_31__I_0_add_566_4 (.CI(n17797), .I0(n838_adj_571[1]), 
            .I1(n108_c), .CO(n17798));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_3_lut (.I0(GND_net), .I1(n835_adj_564[0]), 
            .I2(n105_c), .I3(n17751), .O(n834_adj_574[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_563_15_lut (.I0(GND_net), .I1(n835_adj_564[12]), 
            .I2(n141), .I3(n17763), .O(n834_adj_574[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_8_lut (.I0(GND_net), .I1(n839_adj_570[5]), 
            .I2(n120_c), .I3(n17816), .O(n838_adj_571[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_15 (.CI(n17763), .I0(n835_adj_564[12]), 
            .I1(n141), .CO(n17764));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_14_lut (.I0(GND_net), .I1(n835_adj_564[11]), 
            .I2(n138_c), .I3(n17762), .O(n834_adj_574[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_12 (.CI(n17891), .I0(n843[9]), 
            .I1(n132_c), .CO(n17892));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_11_lut (.I0(GND_net), .I1(n843[8]), 
            .I2(n129_c), .I3(n17890), .O(n842[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_566_3_lut (.I0(GND_net), .I1(n838_adj_571[0]), 
            .I2(n105_c), .I3(n17796), .O(n837_adj_572[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_14 (.CI(n17762), .I0(n835_adj_564[11]), 
            .I1(n138_c), .CO(n17763));
    SB_CARRY Error_sub_temp_31__I_0_add_571_11 (.CI(n17890), .I0(n843[8]), 
            .I1(n129_c), .CO(n17891));
    SB_CARRY Error_sub_temp_31__I_0_add_566_3 (.CI(n17796), .I0(n838_adj_571[0]), 
            .I1(n105_c), .CO(n17797));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_10_lut (.I0(GND_net), .I1(n843[7]), 
            .I2(n126_c), .I3(n17889), .O(n842[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_8 (.CI(n17816), .I0(n839_adj_570[5]), 
            .I1(n120_c), .CO(n17817));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n837_adj_572[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_563_13_lut (.I0(GND_net), .I1(n835_adj_564[10]), 
            .I2(n135_c), .I3(n17761), .O(n834_adj_574[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_10 (.CI(n17889), .I0(n843[7]), 
            .I1(n126_c), .CO(n17890));
    SB_CARRY Error_sub_temp_31__I_0_add_566_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17796));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_9_lut (.I0(GND_net), .I1(n843[6]), 
            .I2(n123_c), .I3(n17888), .O(n842[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_7_lut (.I0(GND_net), .I1(n839_adj_570[4]), 
            .I2(n117_c), .I3(n17815), .O(n838_adj_571[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_9 (.CI(n17888), .I0(n843[6]), 
            .I1(n123_c), .CO(n17889));
    SB_CARRY Error_sub_temp_31__I_0_add_567_7 (.CI(n17815), .I0(n839_adj_570[4]), 
            .I1(n117_c), .CO(n17816));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_8_lut (.I0(GND_net), .I1(n843[5]), 
            .I2(n120_c), .I3(n17887), .O(n842[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_6_lut (.I0(GND_net), .I1(n839_adj_570[3]), 
            .I2(n114_c), .I3(n17814), .O(n838_adj_571[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_8 (.CI(n17541), .I0(n834[5]), 
            .I1(n102_c), .CO(n17542));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_15_lut (.I0(GND_net), .I1(n834[12]), 
            .I2(n102_c), .I3(n17548), .O(n833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_16 (.CI(n17549), .I0(n834[13]), 
            .I1(n741_c), .CO(n743_adj_410));
    SB_CARRY Error_sub_temp_31__I_0_add_571_8 (.CI(n17887), .I0(n843[5]), 
            .I1(n120_c), .CO(n17888));
    SB_CARRY Error_sub_temp_31__I_0_add_567_6 (.CI(n17814), .I0(n839_adj_570[3]), 
            .I1(n114_c), .CO(n17815));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_7_lut (.I0(GND_net), .I1(n835[4]), 
            .I2(n105_c), .I3(n17555), .O(n834[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_13_lut (.I0(GND_net), .I1(n835[10]), 
            .I2(n105_c), .I3(n17561), .O(n834[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_4_lut (.I0(GND_net), .I1(n836[1]), 
            .I2(n108_c), .I3(n17567), .O(n835[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_4 (.CI(n17567), .I0(n836[1]), 
            .I1(n108_c), .CO(n17568));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_7_lut (.I0(GND_net), .I1(n843[4]), 
            .I2(n117_c), .I3(n17886), .O(n842[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_5_lut (.I0(GND_net), .I1(n839_adj_570[2]), 
            .I2(n111_c), .I3(n17813), .O(n838_adj_571[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_15_lut (.I0(GND_net), .I1(n836[12]), 
            .I2(n108_c), .I3(n17578), .O(n835[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_6_lut (.I0(GND_net), .I1(n837[3]), 
            .I2(n111_c), .I3(n17584), .O(n836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_13 (.CI(n17591), .I0(n837[10]), 
            .I1(n111_c), .CO(n17592));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_12_lut (.I0(GND_net), .I1(n837[9]), 
            .I2(n111_c), .I3(n17590), .O(n836[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_7 (.CI(n17886), .I0(n843[4]), 
            .I1(n117_c), .CO(n17887));
    SB_CARRY Error_sub_temp_31__I_0_add_567_5 (.CI(n17813), .I0(n839_adj_570[2]), 
            .I1(n111_c), .CO(n17814));
    SB_CARRY paramCurrentControlP_15__I_0_add_566_13 (.CI(n17606), .I0(n838[10]), 
            .I1(n114_c), .CO(n17607));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_7 (.CI(n17615), .I0(n839[4]), 
            .I1(n117_c), .CO(n17616));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_14 (.CI(n17622), .I0(n839[11]), 
            .I1(n117_c), .CO(n17623));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_13_lut (.I0(GND_net), .I1(n839[10]), 
            .I2(n117_c), .I3(n17621), .O(n838[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_571_6_lut (.I0(GND_net), .I1(n843[3]), 
            .I2(n114_c), .I3(n17885), .O(n842[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_4_lut (.I0(GND_net), .I1(n839_adj_570[1]), 
            .I2(n108_c), .I3(n17812), .O(n838_adj_571[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_9_lut (.I0(GND_net), .I1(n840[6]), 
            .I2(n120_c), .I3(n17632), .O(n839[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_10_lut (.I0(GND_net), .I1(n841[7]), 
            .I2(n123_c), .I3(n17648), .O(n840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_6 (.CI(n17885), .I0(n843[3]), 
            .I1(n114_c), .CO(n17886));
    SB_CARRY Error_sub_temp_31__I_0_add_567_4 (.CI(n17812), .I0(n839_adj_570[1]), 
            .I1(n108_c), .CO(n17813));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_16_lut (.I0(GND_net), .I1(n837_adj_572[13]), 
            .I2(n146), .I3(n17794), .O(n836_adj_565[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_3_lut (.I0(GND_net), .I1(n839_adj_570[0]), 
            .I2(n105_c), .I3(n17811), .O(n838_adj_571[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_571_5_lut (.I0(GND_net), .I1(n843[2]), 
            .I2(n111_c), .I3(n17884), .O(n842[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_5 (.CI(n17884), .I0(n843[2]), 
            .I1(n111_c), .CO(n17885));
    SB_CARRY Error_sub_temp_31__I_0_add_563_3 (.CI(n17751), .I0(n835_adj_564[0]), 
            .I1(n105_c), .CO(n17752));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n834_adj_574[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_571_4_lut (.I0(GND_net), .I1(n843[1]), 
            .I2(n108_c), .I3(n17883), .O(n842[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_3 (.CI(n17811), .I0(n839_adj_570[0]), 
            .I1(n105_c), .CO(n17812));
    SB_CARRY Error_sub_temp_31__I_0_add_565_16 (.CI(n17794), .I0(n837_adj_572[13]), 
            .I1(n146), .CO(n755));
    SB_LUT4 Error_sub_temp_31__I_0_add_567_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n838_adj_571[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_13 (.CI(n17761), .I0(n835_adj_564[10]), 
            .I1(n135_c), .CO(n17762));
    SB_CARRY Error_sub_temp_31__I_0_add_571_4 (.CI(n17883), .I0(n843[1]), 
            .I1(n108_c), .CO(n17884));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_3_lut (.I0(GND_net), .I1(n843[0]), 
            .I2(n105_c), .I3(n17882), .O(n842[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_563_12_lut (.I0(GND_net), .I1(n835_adj_564[9]), 
            .I2(n132_c), .I3(n17760), .O(n834_adj_574[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_15_lut (.I0(GND_net), .I1(n837_adj_572[12]), 
            .I2(n141), .I3(n17793), .O(n836_adj_565[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_567_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17811));
    SB_LUT4 Error_sub_temp_31__I_0_add_566_16_lut (.I0(GND_net), .I1(n838_adj_571[13]), 
            .I2(n146), .I3(n17809), .O(n837_adj_572[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_3 (.CI(n17882), .I0(n843[0]), 
            .I1(n105_c), .CO(n17883));
    SB_LUT4 Error_sub_temp_31__I_0_add_571_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n842[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_571_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17882));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_6 (.CI(n17584), .I0(n837[3]), 
            .I1(n111_c), .CO(n17585));
    SB_CARRY Error_sub_temp_31__I_0_add_566_16 (.CI(n17809), .I0(n838_adj_571[13]), 
            .I1(n146), .CO(n759_adj_354));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_12 (.CI(n17590), .I0(n837[9]), 
            .I1(n111_c), .CO(n17591));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_12_lut (.I0(GND_net), .I1(n838[9]), 
            .I2(n114_c), .I3(n17605), .O(n837[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_570_16_lut (.I0(GND_net), .I1(n842[13]), 
            .I2(n146), .I3(n17880), .O(n841_adj_568[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_15 (.CI(n17793), .I0(n837_adj_572[12]), 
            .I1(n141), .CO(n17794));
    SB_CARRY Error_sub_temp_31__I_0_add_570_16 (.CI(n17880), .I0(n842[13]), 
            .I1(n146), .CO(n775));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_15_lut (.I0(GND_net), .I1(n842[12]), 
            .I2(n141), .I3(n17879), .O(n841_adj_568[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_15 (.CI(n17879), .I0(n842[12]), 
            .I1(n141), .CO(n17880));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_14_lut (.I0(GND_net), .I1(n842[11]), 
            .I2(n138_c), .I3(n17878), .O(n841_adj_568[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_14 (.CI(n17878), .I0(n842[11]), 
            .I1(n138_c), .CO(n17879));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_13_lut (.I0(GND_net), .I1(n842[10]), 
            .I2(n135_c), .I3(n17877), .O(n841_adj_568[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_13 (.CI(n17877), .I0(n842[10]), 
            .I1(n135_c), .CO(n17878));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_12_lut (.I0(GND_net), .I1(n842[9]), 
            .I2(n132_c), .I3(n17876), .O(n841_adj_568[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_12 (.CI(n17876), .I0(n842[9]), 
            .I1(n132_c), .CO(n17877));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_11_lut (.I0(GND_net), .I1(n842[8]), 
            .I2(n129_c), .I3(n17875), .O(n841_adj_568[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_566_13_lut (.I0(GND_net), .I1(n838_adj_571[10]), 
            .I2(n135_c), .I3(n17806), .O(n837_adj_572[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_11 (.CI(n17875), .I0(n842[8]), 
            .I1(n129_c), .CO(n17876));
    SB_CARRY Error_sub_temp_31__I_0_add_566_14 (.CI(n17807), .I0(n838_adj_571[11]), 
            .I1(n138_c), .CO(n17808));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_10_lut (.I0(GND_net), .I1(n842[7]), 
            .I2(n126_c), .I3(n17874), .O(n841_adj_568[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_566_14_lut (.I0(GND_net), .I1(n838_adj_571[11]), 
            .I2(n138_c), .I3(n17807), .O(n837_adj_572[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_566_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_7_lut (.I0(GND_net), .I1(n834[4]), 
            .I2(n102_c), .I3(n17540), .O(n833[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_16_lut (.I0(GND_net), .I1(n834[13]), 
            .I2(n741_c), .I3(n17549), .O(n833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_7 (.CI(n17555), .I0(n835[4]), 
            .I1(n105_c), .CO(n17556));
    SB_CARRY Error_sub_temp_31__I_0_add_570_10 (.CI(n17874), .I0(n842[7]), 
            .I1(n126_c), .CO(n17875));
    SB_CARRY Error_sub_temp_31__I_0_add_563_12 (.CI(n17760), .I0(n835_adj_564[9]), 
            .I1(n132_c), .CO(n17761));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_6_lut (.I0(GND_net), .I1(n835[3]), 
            .I2(n105_c), .I3(n17554), .O(n834[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_13 (.CI(n17561), .I0(n835[10]), 
            .I1(n105_c), .CO(n17562));
    SB_CARRY paramCurrentControlP_15__I_0_add_564_15 (.CI(n17578), .I0(n836[12]), 
            .I1(n108_c), .CO(n17579));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_3_lut (.I0(GND_net), .I1(n836[0]), 
            .I2(n108_c), .I3(n17566), .O(n835[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_570_9_lut (.I0(GND_net), .I1(n842[6]), 
            .I2(n123_c), .I3(n17873), .O(n841_adj_568[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_566_15 (.CI(n17808), .I0(n838_adj_571[12]), 
            .I1(n141), .CO(n17809));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_14_lut (.I0(GND_net), .I1(n836[11]), 
            .I2(n108_c), .I3(n17577), .O(n835[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_5_lut (.I0(GND_net), .I1(n837[2]), 
            .I2(n111_c), .I3(n17583), .O(n836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_12 (.CI(n17605), .I0(n838[9]), 
            .I1(n114_c), .CO(n17606));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_11_lut (.I0(GND_net), .I1(n837[8]), 
            .I2(n111_c), .I3(n17589), .O(n836[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_9 (.CI(n17873), .I0(n842[6]), 
            .I1(n123_c), .CO(n17874));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_11_lut (.I0(GND_net), .I1(n835_adj_564[8]), 
            .I2(n129_c), .I3(n17759), .O(n834_adj_574[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_11_lut (.I0(GND_net), .I1(n838[8]), 
            .I2(n114_c), .I3(n17604), .O(n837[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_6_lut (.I0(GND_net), .I1(n839[3]), 
            .I2(n117_c), .I3(n17614), .O(n838[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_9 (.CI(n17632), .I0(n840[6]), 
            .I1(n120_c), .CO(n17633));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_13 (.CI(n17621), .I0(n839[10]), 
            .I1(n117_c), .CO(n17622));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_8_lut (.I0(GND_net), .I1(n842[5]), 
            .I2(n120_c), .I3(n17872), .O(n841_adj_568[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_14_lut (.I0(GND_net), .I1(n837_adj_572[11]), 
            .I2(n138_c), .I3(n17792), .O(n836_adj_565[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_10 (.CI(n17648), .I0(n841[7]), 
            .I1(n123_c), .CO(n17649));
    SB_CARRY Error_sub_temp_31__I_0_add_570_8 (.CI(n17872), .I0(n842[5]), 
            .I1(n120_c), .CO(n17873));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_7_lut (.I0(GND_net), .I1(n842[4]), 
            .I2(n117_c), .I3(n17871), .O(n841_adj_568[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_8_lut (.I0(GND_net), .I1(n840[5]), 
            .I2(n120_c), .I3(n17631), .O(n839[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_9_lut (.I0(GND_net), .I1(n841[6]), 
            .I2(n123_c), .I3(n17647), .O(n840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_7 (.CI(n17871), .I0(n842[4]), 
            .I1(n117_c), .CO(n17872));
    SB_CARRY Error_sub_temp_31__I_0_add_565_14 (.CI(n17792), .I0(n837_adj_572[11]), 
            .I1(n138_c), .CO(n17793));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_6_lut (.I0(GND_net), .I1(n842[3]), 
            .I2(n114_c), .I3(n17870), .O(n841_adj_568[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_6 (.CI(n17870), .I0(n842[3]), 
            .I1(n114_c), .CO(n17871));
    SB_CARRY Error_sub_temp_31__I_0_add_563_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17751));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_13_lut (.I0(GND_net), .I1(n837_adj_572[10]), 
            .I2(n135_c), .I3(n17791), .O(n836_adj_565[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_11 (.CI(n17759), .I0(n835_adj_564[8]), 
            .I1(n129_c), .CO(n17760));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_5_lut (.I0(GND_net), .I1(n842[2]), 
            .I2(n111_c), .I3(n17869), .O(n841_adj_568[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_9 (.CI(n17647), .I0(n841[6]), 
            .I1(n123_c), .CO(n17648));
    SB_CARRY Error_sub_temp_31__I_0_add_570_5 (.CI(n17869), .I0(n842[2]), 
            .I1(n111_c), .CO(n17870));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_4_lut (.I0(GND_net), .I1(n842[1]), 
            .I2(n108_c), .I3(n17868), .O(n841_adj_568[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_4 (.CI(n17868), .I0(n842[1]), 
            .I1(n108_c), .CO(n17869));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_3_lut (.I0(GND_net), .I1(n842[0]), 
            .I2(n105_c), .I3(n17867), .O(n841_adj_568[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_11 (.CI(n17604), .I0(n838[8]), 
            .I1(n114_c), .CO(n17605));
    SB_CARRY paramCurrentControlP_15__I_0_add_568_8 (.CI(n17631), .I0(n840[5]), 
            .I1(n120_c), .CO(n17632));
    SB_CARRY Error_sub_temp_31__I_0_add_570_3 (.CI(n17867), .I0(n842[0]), 
            .I1(n105_c), .CO(n17868));
    SB_LUT4 Error_sub_temp_31__I_0_add_570_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n841_adj_568[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_570_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17867));
    SB_CARRY Error_sub_temp_31__I_0_add_565_13 (.CI(n17791), .I0(n837_adj_572[10]), 
            .I1(n135_c), .CO(n17792));
    SB_DFF currentControlITerm_i6 (.Q(currentControlITerm[6]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14325));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_DFF currentControlITerm_i0 (.Q(currentControlITerm[0]), .C(pin3_clk_16mhz_N_keep), 
           .D(n19782));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_LUT4 paramCurrentControlP_15__I_0_i522_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[24]), .I2(GND_net), .I3(GND_net), .O(n769_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i522_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_547_27_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[25]), 
            .I2(currentControlITerm[31]), .I3(n15592), .O(preSatVoltage[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_28 (.CI(n15593), .I0(Proportional_Gain_mul_temp[26]), 
            .I1(currentControlITerm[31]), .CO(n15594));
    SB_LUT4 add_547_28_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[26]), 
            .I2(currentControlITerm[31]), .I3(n15593), .O(preSatVoltage[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_29 (.CI(n15594), .I0(Proportional_Gain_mul_temp[27]), 
            .I1(currentControlITerm[31]), .CO(n15595));
    SB_LUT4 add_547_29_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[27]), 
            .I2(currentControlITerm[31]), .I3(n15594), .O(preSatVoltage[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_30 (.CI(n15595), .I0(Proportional_Gain_mul_temp[28]), 
            .I1(currentControlITerm[31]), .CO(n15596));
    SB_LUT4 add_547_30_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[28]), 
            .I2(currentControlITerm[31]), .I3(n15595), .O(preSatVoltage[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_547_31_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[29]), 
            .I2(currentControlITerm[31]), .I3(n15596), .O(preSatVoltage[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_547_31 (.CI(n15596), .I0(Proportional_Gain_mul_temp[29]), 
            .I1(currentControlITerm[31]), .CO(n15597));
    SB_DFF currentControlITerm_i5 (.Q(currentControlITerm[5]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14324));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_CARRY paramCurrentControlP_15__I_0_add_562_7 (.CI(n17540), .I0(n834[4]), 
            .I1(n102_c), .CO(n17541));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_6_lut (.I0(GND_net), .I1(n834[3]), 
            .I2(n102_c), .I3(n17539), .O(n833[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_2 (.CI(GND_net), .I0(n108_c), 
            .I1(n105_c), .CO(n17551));
    SB_CARRY paramCurrentControlP_15__I_0_add_563_6 (.CI(n17554), .I0(n835[3]), 
            .I1(n105_c), .CO(n17555));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_12_lut (.I0(GND_net), .I1(n835[9]), 
            .I2(n105_c), .I3(n17560), .O(n834[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_6 (.CI(n17614), .I0(n839[3]), 
            .I1(n117_c), .CO(n17615));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_10_lut (.I0(GND_net), .I1(n838[7]), 
            .I2(n114_c), .I3(n17603), .O(n837[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_10 (.CI(n17603), .I0(n838[7]), 
            .I1(n114_c), .CO(n17604));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_9_lut (.I0(GND_net), .I1(n838[6]), 
            .I2(n114_c), .I3(n17602), .O(n837[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_9 (.CI(n17602), .I0(n838[6]), 
            .I1(n114_c), .CO(n17603));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_8_lut (.I0(GND_net), .I1(n838[5]), 
            .I2(n114_c), .I3(n17601), .O(n837[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_8 (.CI(n17601), .I0(n838[5]), 
            .I1(n114_c), .CO(n17602));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_7_lut (.I0(GND_net), .I1(n838[4]), 
            .I2(n114_c), .I3(n17600), .O(n837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_7 (.CI(n17600), .I0(n838[4]), 
            .I1(n114_c), .CO(n17601));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_6_lut (.I0(GND_net), .I1(n838[3]), 
            .I2(n114_c), .I3(n17599), .O(n837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_6 (.CI(n17599), .I0(n838[3]), 
            .I1(n114_c), .CO(n17600));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_5_lut (.I0(GND_net), .I1(n838[2]), 
            .I2(n114_c), .I3(n17598), .O(n837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_5 (.CI(n17598), .I0(n838[2]), 
            .I1(n114_c), .CO(n17599));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_4_lut (.I0(GND_net), .I1(n838[1]), 
            .I2(n114_c), .I3(n17597), .O(n837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_4 (.CI(n17597), .I0(n838[1]), 
            .I1(n114_c), .CO(n17598));
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_3_lut (.I0(GND_net), .I1(n838[0]), 
            .I2(n114_c), .I3(n17596), .O(n837[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_12 (.CI(n17560), .I0(n835[9]), 
            .I1(n105_c), .CO(n17561));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_8_lut (.I0(GND_net), .I1(n841[5]), 
            .I2(n123_c), .I3(n17646), .O(n840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_3 (.CI(n17566), .I0(n836[0]), 
            .I1(n108_c), .CO(n17567));
    SB_CARRY paramCurrentControlP_15__I_0_add_564_14 (.CI(n17577), .I0(n836[11]), 
            .I1(n108_c), .CO(n17578));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_5 (.CI(n17583), .I0(n837[2]), 
            .I1(n111_c), .CO(n17584));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_4_lut (.I0(GND_net), .I1(n837[1]), 
            .I2(n111_c), .I3(n17582), .O(n836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_7_lut (.I0(GND_net), .I1(n840[4]), 
            .I2(n120_c), .I3(n17630), .O(n839[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_11 (.CI(n17589), .I0(n837[8]), 
            .I1(n111_c), .CO(n17590));
    SB_CARRY paramCurrentControlP_15__I_0_add_566_3 (.CI(n17596), .I0(n838[0]), 
            .I1(n114_c), .CO(n17597));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_5_lut (.I0(GND_net), .I1(n839[2]), 
            .I2(n117_c), .I3(n17613), .O(n838[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_5 (.CI(n17613), .I0(n839[2]), 
            .I1(n117_c), .CO(n17614));
    SB_CARRY paramCurrentControlP_15__I_0_add_562_6 (.CI(n17539), .I0(n834[3]), 
            .I1(n102_c), .CO(n17540));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_12_lut (.I0(GND_net), .I1(n837_adj_572[9]), 
            .I2(n132_c), .I3(n17790), .O(n836_adj_565[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_2_lut (.I0(GND_net), .I1(n108_c), 
            .I2(n105_c), .I3(GND_net), .O(n834[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_12_lut (.I0(GND_net), .I1(n839[9]), 
            .I2(n117_c), .I3(n17620), .O(n838[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_12 (.CI(n17620), .I0(n839[9]), 
            .I1(n117_c), .CO(n17621));
    SB_CARRY paramCurrentControlP_15__I_0_add_568_7 (.CI(n17630), .I0(n840[4]), 
            .I1(n120_c), .CO(n17631));
    SB_CARRY paramCurrentControlP_15__I_0_add_569_8 (.CI(n17646), .I0(n841[5]), 
            .I1(n123_c), .CO(n17647));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_11_lut (.I0(GND_net), .I1(n834[8]), 
            .I2(n102_c), .I3(n17544), .O(n833[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_12 (.CI(n17790), .I0(n837_adj_572[9]), 
            .I1(n132_c), .CO(n17791));
    SB_CARRY paramCurrentControlP_15__I_0_add_562_11 (.CI(n17544), .I0(n834[8]), 
            .I1(n102_c), .CO(n17545));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_16_lut (.I0(GND_net), .I1(n834_adj_574[13]), 
            .I2(n146), .I3(n17749), .O(n833_adj_575[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_16 (.CI(n17749), .I0(n834_adj_574[13]), 
            .I1(n146), .CO(n743));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_7_lut (.I0(GND_net), .I1(n841[4]), 
            .I2(n123_c), .I3(n17645), .O(n840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_563_10_lut (.I0(GND_net), .I1(n835_adj_564[7]), 
            .I2(n126_c), .I3(n17758), .O(n834_adj_574[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_11_lut (.I0(GND_net), .I1(n837_adj_572[8]), 
            .I2(n129_c), .I3(n17789), .O(n836_adj_565[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_6_lut (.I0(GND_net), .I1(n840[3]), 
            .I2(n120_c), .I3(n17629), .O(n839[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_11_lut (.I0(GND_net), .I1(n835[8]), 
            .I2(n105_c), .I3(n17559), .O(n834[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_11_lut (.I0(GND_net), .I1(n839[8]), 
            .I2(n117_c), .I3(n17619), .O(n838[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_569_16_lut (.I0(GND_net), .I1(n841_adj_568[13]), 
            .I2(n146), .I3(n17854), .O(n840_adj_569[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_16 (.CI(n17854), .I0(n841_adj_568[13]), 
            .I1(n146), .CO(n771_adj_353));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_15_lut (.I0(GND_net), .I1(n841_adj_568[12]), 
            .I2(n141), .I3(n17853), .O(n840_adj_569[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_15 (.CI(n17853), .I0(n841_adj_568[12]), 
            .I1(n141), .CO(n17854));
    SB_CARRY paramCurrentControlP_15__I_0_add_568_6 (.CI(n17629), .I0(n840[3]), 
            .I1(n120_c), .CO(n17630));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_14_lut (.I0(GND_net), .I1(n841_adj_568[11]), 
            .I2(n138_c), .I3(n17852), .O(n840_adj_569[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_5_lut (.I0(GND_net), .I1(n840[2]), 
            .I2(n120_c), .I3(n17628), .O(n839[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_14 (.CI(n17852), .I0(n841_adj_568[11]), 
            .I1(n138_c), .CO(n17853));
    SB_CARRY Error_sub_temp_31__I_0_add_565_11 (.CI(n17789), .I0(n837_adj_572[8]), 
            .I1(n129_c), .CO(n17790));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_2_lut (.I0(GND_net), .I1(n111_c), 
            .I2(n108_c), .I3(GND_net), .O(n835[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_7 (.CI(n17645), .I0(n841[4]), 
            .I1(n123_c), .CO(n17646));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_13_lut (.I0(GND_net), .I1(n841_adj_568[10]), 
            .I2(n135_c), .I3(n17851), .O(n840_adj_569[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_13 (.CI(n17851), .I0(n841_adj_568[10]), 
            .I1(n135_c), .CO(n17852));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_12_lut (.I0(GND_net), .I1(n841_adj_568[9]), 
            .I2(n132_c), .I3(n17850), .O(n840_adj_569[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_12 (.CI(n17850), .I0(n841_adj_568[9]), 
            .I1(n132_c), .CO(n17851));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_11_lut (.I0(GND_net), .I1(n841_adj_568[8]), 
            .I2(n129_c), .I3(n17849), .O(n840_adj_569[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_11 (.CI(n17849), .I0(n841_adj_568[8]), 
            .I1(n129_c), .CO(n17850));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_10_lut (.I0(GND_net), .I1(n841_adj_568[7]), 
            .I2(n126_c), .I3(n17848), .O(n840_adj_569[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_10 (.CI(n17848), .I0(n841_adj_568[7]), 
            .I1(n126_c), .CO(n17849));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_9_lut (.I0(GND_net), .I1(n841_adj_568[6]), 
            .I2(n123_c), .I3(n17847), .O(n840_adj_569[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_9 (.CI(n17847), .I0(n841_adj_568[6]), 
            .I1(n123_c), .CO(n17848));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_8_lut (.I0(GND_net), .I1(n841_adj_568[5]), 
            .I2(n120_c), .I3(n17846), .O(n840_adj_569[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_8 (.CI(n17846), .I0(n841_adj_568[5]), 
            .I1(n120_c), .CO(n17847));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_13_lut (.I0(GND_net), .I1(n836[10]), 
            .I2(n108_c), .I3(n17576), .O(n835[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_569_7_lut (.I0(GND_net), .I1(n841_adj_568[4]), 
            .I2(n117_c), .I3(n17845), .O(n840_adj_569[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_13 (.CI(n17576), .I0(n836[10]), 
            .I1(n108_c), .CO(n17577));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_5_lut (.I0(GND_net), .I1(n834[2]), 
            .I2(n102_c), .I3(n17538), .O(n833[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_3 (.CI(n17551), .I0(n835[0]), 
            .I1(n105_c), .CO(n17552));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_10_lut (.I0(GND_net), .I1(n834[7]), 
            .I2(n102_c), .I3(n17543), .O(n833[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_10 (.CI(n17543), .I0(n834[7]), 
            .I1(n102_c), .CO(n17544));
    SB_CARRY Error_sub_temp_31__I_0_add_569_7 (.CI(n17845), .I0(n841_adj_568[4]), 
            .I1(n117_c), .CO(n17846));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_6_lut (.I0(GND_net), .I1(n841[3]), 
            .I2(n123_c), .I3(n17644), .O(n840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_563_11 (.CI(n17559), .I0(n835[8]), 
            .I1(n105_c), .CO(n17560));
    SB_CARRY paramCurrentControlP_15__I_0_add_564_2 (.CI(GND_net), .I0(n111_c), 
            .I1(n108_c), .CO(n17566));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_12_lut (.I0(GND_net), .I1(n836[9]), 
            .I2(n108_c), .I3(n17575), .O(n835[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_564_12 (.CI(n17575), .I0(n836[9]), 
            .I1(n108_c), .CO(n17576));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_6_lut (.I0(GND_net), .I1(n841_adj_568[3]), 
            .I2(n114_c), .I3(n17844), .O(n840_adj_569[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_5 (.CI(n17628), .I0(n840[2]), 
            .I1(n120_c), .CO(n17629));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_4 (.CI(n17582), .I0(n837[1]), 
            .I1(n111_c), .CO(n17583));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_10_lut (.I0(GND_net), .I1(n837[7]), 
            .I2(n111_c), .I3(n17588), .O(n836[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_2_lut (.I0(GND_net), .I1(n117_c), 
            .I2(n114_c), .I3(GND_net), .O(n837[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_566_2 (.CI(GND_net), .I0(n117_c), 
            .I1(n114_c), .CO(n17596));
    SB_CARRY Error_sub_temp_31__I_0_add_569_6 (.CI(n17844), .I0(n841_adj_568[3]), 
            .I1(n114_c), .CO(n17845));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_3_lut (.I0(GND_net), .I1(n837[0]), 
            .I2(n111_c), .I3(n17581), .O(n836[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_10_lut (.I0(GND_net), .I1(n837_adj_572[7]), 
            .I2(n126_c), .I3(n17788), .O(n836_adj_565[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_10 (.CI(n17588), .I0(n837[7]), 
            .I1(n111_c), .CO(n17589));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_4_lut (.I0(GND_net), .I1(n839[1]), 
            .I2(n117_c), .I3(n17612), .O(n838[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_569_5_lut (.I0(GND_net), .I1(n841_adj_568[2]), 
            .I2(n111_c), .I3(n17843), .O(n840_adj_569[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_5 (.CI(n17843), .I0(n841_adj_568[2]), 
            .I1(n111_c), .CO(n17844));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_4 (.CI(n17612), .I0(n839[1]), 
            .I1(n117_c), .CO(n17613));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_11 (.CI(n17619), .I0(n839[8]), 
            .I1(n117_c), .CO(n17620));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_4_lut (.I0(GND_net), .I1(n840[1]), 
            .I2(n120_c), .I3(n17627), .O(n839[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_6 (.CI(n17644), .I0(n841[3]), 
            .I1(n123_c), .CO(n17645));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_5_lut (.I0(GND_net), .I1(n841[2]), 
            .I2(n123_c), .I3(n17643), .O(n840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_569_4_lut (.I0(GND_net), .I1(n841_adj_568[1]), 
            .I2(n108_c), .I3(n17842), .O(n840_adj_569[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_16_lut (.I0(GND_net), .I1(n837[13]), 
            .I2(n753_c), .I3(n17594), .O(n836[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_10 (.CI(n17788), .I0(n837_adj_572[7]), 
            .I1(n126_c), .CO(n17789));
    SB_CARRY paramCurrentControlP_15__I_0_add_565_16 (.CI(n17594), .I0(n837[13]), 
            .I1(n753_c), .CO(n755_adj_404));
    SB_CARRY Error_sub_temp_31__I_0_add_569_4 (.CI(n17842), .I0(n841_adj_568[1]), 
            .I1(n108_c), .CO(n17843));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_3_lut (.I0(GND_net), .I1(n841_adj_568[0]), 
            .I2(n105_c), .I3(n17841), .O(n840_adj_569[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_3 (.CI(n17841), .I0(n841_adj_568[0]), 
            .I1(n105_c), .CO(n17842));
    SB_CARRY paramCurrentControlP_15__I_0_add_569_5 (.CI(n17643), .I0(n841[2]), 
            .I1(n123_c), .CO(n17644));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_15_lut (.I0(GND_net), .I1(n834_adj_574[12]), 
            .I2(n141), .I3(n17748), .O(n833_adj_575[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_10 (.CI(n17758), .I0(n835_adj_564[7]), 
            .I1(n126_c), .CO(n17759));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_9_lut (.I0(GND_net), .I1(n837_adj_572[6]), 
            .I2(n123_c), .I3(n17787), .O(n836_adj_565[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_9 (.CI(n17787), .I0(n837_adj_572[6]), 
            .I1(n123_c), .CO(n17788));
    SB_LUT4 Error_sub_temp_31__I_0_add_569_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n840_adj_569[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_569_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17841));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_16_lut (.I0(GND_net), .I1(n840_adj_569[13]), 
            .I2(n146), .I3(n17839), .O(n839_adj_570[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_4 (.CI(n17627), .I0(n840[1]), 
            .I1(n120_c), .CO(n17628));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_4_lut (.I0(GND_net), .I1(n841[1]), 
            .I2(n123_c), .I3(n17642), .O(n840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_16 (.CI(n17839), .I0(n840_adj_569[13]), 
            .I1(n146), .CO(n767));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_15_lut (.I0(GND_net), .I1(n840_adj_569[12]), 
            .I2(n141), .I3(n17838), .O(n839_adj_570[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_15 (.CI(n17838), .I0(n840_adj_569[12]), 
            .I1(n141), .CO(n17839));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_14_lut (.I0(GND_net), .I1(n840_adj_569[11]), 
            .I2(n138_c), .I3(n17837), .O(n839_adj_570[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_14 (.CI(n17837), .I0(n840_adj_569[11]), 
            .I1(n138_c), .CO(n17838));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_13_lut (.I0(GND_net), .I1(n840_adj_569[10]), 
            .I2(n135_c), .I3(n17836), .O(n839_adj_570[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_13 (.CI(n17836), .I0(n840_adj_569[10]), 
            .I1(n135_c), .CO(n17837));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_12_lut (.I0(GND_net), .I1(n840_adj_569[9]), 
            .I2(n132_c), .I3(n17835), .O(n839_adj_570[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_12 (.CI(n17835), .I0(n840_adj_569[9]), 
            .I1(n132_c), .CO(n17836));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_11_lut (.I0(GND_net), .I1(n840_adj_569[8]), 
            .I2(n129_c), .I3(n17834), .O(n839_adj_570[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_11 (.CI(n17834), .I0(n840_adj_569[8]), 
            .I1(n129_c), .CO(n17835));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_10_lut (.I0(GND_net), .I1(n840_adj_569[7]), 
            .I2(n126_c), .I3(n17833), .O(n839_adj_570[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_10 (.CI(n17833), .I0(n840_adj_569[7]), 
            .I1(n126_c), .CO(n17834));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_9_lut (.I0(GND_net), .I1(n840_adj_569[6]), 
            .I2(n123_c), .I3(n17832), .O(n839_adj_570[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_9 (.CI(n17832), .I0(n840_adj_569[6]), 
            .I1(n123_c), .CO(n17833));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_8_lut (.I0(GND_net), .I1(n840_adj_569[5]), 
            .I2(n120_c), .I3(n17831), .O(n839_adj_570[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_8_lut (.I0(GND_net), .I1(n837_adj_572[5]), 
            .I2(n120_c), .I3(n17786), .O(n836_adj_565[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_3_lut (.I0(GND_net), .I1(n839[0]), 
            .I2(n117_c), .I3(n17611), .O(n838[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_5 (.CI(n17538), .I0(n834[2]), 
            .I1(n102_c), .CO(n17539));
    SB_CARRY Error_sub_temp_31__I_0_add_568_8 (.CI(n17831), .I0(n840_adj_569[5]), 
            .I1(n120_c), .CO(n17832));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_7_lut (.I0(GND_net), .I1(n840_adj_569[4]), 
            .I2(n117_c), .I3(n17830), .O(n839_adj_570[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_4_lut (.I0(GND_net), .I1(n834[1]), 
            .I2(n102_c), .I3(n17537), .O(n833[2])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_4 (.CI(n17537), .I0(n834[1]), 
            .I1(n102_c), .CO(n17538));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_9_lut (.I0(GND_net), .I1(n834[6]), 
            .I2(n102_c), .I3(n17542), .O(n833[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_10_lut (.I0(GND_net), .I1(n835[7]), 
            .I2(n105_c), .I3(n17558), .O(n834[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_7 (.CI(n17830), .I0(n840_adj_569[4]), 
            .I1(n117_c), .CO(n17831));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_3 (.CI(n17611), .I0(n839[0]), 
            .I1(n117_c), .CO(n17612));
    SB_CARRY Error_sub_temp_31__I_0_add_565_8 (.CI(n17786), .I0(n837_adj_572[5]), 
            .I1(n120_c), .CO(n17787));
    SB_CARRY paramCurrentControlP_15__I_0_add_569_4 (.CI(n17642), .I0(n841[1]), 
            .I1(n123_c), .CO(n17643));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_16_lut (.I0(GND_net), .I1(n835[13]), 
            .I2(n745_c), .I3(n17564), .O(n834[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_568_6_lut (.I0(GND_net), .I1(n840_adj_569[3]), 
            .I2(n114_c), .I3(n17829), .O(n839_adj_570[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_6 (.CI(n17829), .I0(n840_adj_569[3]), 
            .I1(n114_c), .CO(n17830));
    SB_CARRY paramCurrentControlP_15__I_0_add_563_16 (.CI(n17564), .I0(n835[13]), 
            .I1(n745_c), .CO(n747_adj_408));
    SB_LUT4 paramCurrentControlP_15__I_0_add_564_11_lut (.I0(GND_net), .I1(n836[8]), 
            .I2(n108_c), .I3(n17574), .O(n835[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_564_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_9_lut (.I0(GND_net), .I1(n837[6]), 
            .I2(n111_c), .I3(n17587), .O(n836[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_568_5_lut (.I0(GND_net), .I1(n840_adj_569[2]), 
            .I2(n111_c), .I3(n17828), .O(n839_adj_570[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_10_lut (.I0(GND_net), .I1(n839[7]), 
            .I2(n117_c), .I3(n17618), .O(n838[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_565_9 (.CI(n17587), .I0(n837[6]), 
            .I1(n111_c), .CO(n17588));
    SB_LUT4 paramCurrentControlP_15__I_0_add_565_15_lut (.I0(GND_net), .I1(n837[12]), 
            .I2(n111_c), .I3(n17593), .O(n836[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_565_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_567_10 (.CI(n17618), .I0(n839[7]), 
            .I1(n117_c), .CO(n17619));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_2_lut (.I0(GND_net), .I1(n120_c), 
            .I2(n117_c), .I3(GND_net), .O(n838[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_5 (.CI(n17828), .I0(n840_adj_569[2]), 
            .I1(n111_c), .CO(n17829));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n837_adj_572[4]), 
            .I2(n117_c), .I3(n17785), .O(n836_adj_565[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_3_lut (.I0(GND_net), .I1(n840[0]), 
            .I2(n120_c), .I3(n17626), .O(n839[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_3 (.CI(n17626), .I0(n840[0]), 
            .I1(n120_c), .CO(n17627));
    SB_LUT4 Error_sub_temp_31__I_0_add_568_4_lut (.I0(GND_net), .I1(n840_adj_569[1]), 
            .I2(n108_c), .I3(n17827), .O(n839_adj_570[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17826));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_2_lut (.I0(GND_net), .I1(n123_c), 
            .I2(n120_c), .I3(GND_net), .O(n839[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_565_7 (.CI(n17785), .I0(n837_adj_572[4]), 
            .I1(n117_c), .CO(n17786));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_2 (.CI(GND_net), .I0(n120_c), 
            .I1(n117_c), .CO(n17611));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_3_lut (.I0(GND_net), .I1(n841[0]), 
            .I2(n123_c), .I3(n17641), .O(n840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_568_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n839_adj_570[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_3 (.CI(n17826), .I0(n840_adj_569[0]), 
            .I1(n105_c), .CO(n17827));
    SB_CARRY paramCurrentControlP_15__I_0_add_569_3 (.CI(n17641), .I0(n841[0]), 
            .I1(n123_c), .CO(n17642));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n837_adj_572[3]), 
            .I2(n114_c), .I3(n17784), .O(n836_adj_565[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_15 (.CI(n17748), .I0(n834_adj_574[12]), 
            .I1(n141), .CO(n17749));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_14_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[11]), .I2(n138_c), .I3(n17747), .O(Switch_out1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_565_6 (.CI(n17784), .I0(n837_adj_572[3]), 
            .I1(n114_c), .CO(n17785));
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_2_lut (.I0(GND_net), .I1(n126_c), 
            .I2(n123_c), .I3(GND_net), .O(n840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_14 (.CI(n17747), .I0(n834_adj_574[11]), 
            .I1(n138_c), .CO(n17748));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_9_lut (.I0(GND_net), .I1(n835_adj_564[6]), 
            .I2(n123_c), .I3(n17757), .O(n834_adj_574[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n837_adj_572[2]), 
            .I2(n111_c), .I3(n17783), .O(n836_adj_565[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_9_lut (.I0(GND_net), .I1(n839[6]), 
            .I2(n117_c), .I3(n17617), .O(n838[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_9 (.CI(n17757), .I0(n835_adj_564[6]), 
            .I1(n123_c), .CO(n17758));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_8_lut (.I0(GND_net), .I1(n835_adj_564[5]), 
            .I2(n120_c), .I3(n17756), .O(n834_adj_574[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_562_13_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[10]), .I2(n135_c), .I3(n17746), .O(Switch_out1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_563_6 (.CI(n17754), .I0(n835_adj_564[3]), 
            .I1(n114_c), .CO(n17755));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_6_lut (.I0(GND_net), .I1(n835_adj_564[3]), 
            .I2(n114_c), .I3(n17754), .O(n834_adj_574[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_567_16_lut (.I0(GND_net), .I1(n839_adj_570[13]), 
            .I2(n146), .I3(n17824), .O(n838_adj_571[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_2 (.CI(GND_net), .I0(n123_c), 
            .I1(n120_c), .CO(n17626));
    SB_CARRY Error_sub_temp_31__I_0_add_565_5 (.CI(n17783), .I0(n837_adj_572[2]), 
            .I1(n111_c), .CO(n17784));
    SB_LUT4 paramCurrentControlP_15__I_0_add_567_16_lut (.I0(GND_net), .I1(n839[13]), 
            .I2(n761_c), .I3(n17624), .O(n838[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_567_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_563_7 (.CI(n17755), .I0(n835_adj_564[4]), 
            .I1(n117_c), .CO(n17756));
    SB_CARRY Error_sub_temp_31__I_0_add_562_13 (.CI(n17746), .I0(n834_adj_574[10]), 
            .I1(n135_c), .CO(n17747));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_12_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[9]), .I2(n132_c), .I3(n17745), .O(Switch_out1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_12 (.CI(n17745), .I0(n834_adj_574[9]), 
            .I1(n132_c), .CO(n17746));
    SB_LUT4 Error_sub_temp_31__I_0_add_563_7_lut (.I0(GND_net), .I1(n835_adj_564[4]), 
            .I2(n117_c), .I3(n17755), .O(n834_adj_574[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_562_11_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[8]), .I2(n129_c), .I3(n17744), .O(Switch_out1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY paramCurrentControlP_15__I_0_add_569_2 (.CI(GND_net), .I0(n126_c), 
            .I1(n123_c), .CO(n17641));
    SB_LUT4 Error_sub_temp_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n837_adj_572[1]), 
            .I2(n108_c), .I3(n17782), .O(n836_adj_565[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_568_3_lut (.I0(GND_net), .I1(n840_adj_569[0]), 
            .I2(n105_c), .I3(n17826), .O(n839_adj_570[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_568_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_568_4 (.CI(n17827), .I0(n840_adj_569[1]), 
            .I1(n108_c), .CO(n17828));
    SB_CARRY Error_sub_temp_31__I_0_add_562_11 (.CI(n17744), .I0(n834_adj_574[8]), 
            .I1(n129_c), .CO(n17745));
    SB_CARRY Error_sub_temp_31__I_0_add_565_4 (.CI(n17782), .I0(n837_adj_572[1]), 
            .I1(n108_c), .CO(n17783));
    SB_LUT4 add_4257_17_lut (.I0(Not_Equal_relop1_N_201), .I1(n796), .I2(n795), 
            .I3(n17726), .O(Switch_out1[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Error_sub_temp_31__I_0_add_562_10_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[7]), .I2(n126_c), .I3(n17743), .O(Switch_out1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n837_adj_572[0]), 
            .I2(n105_c), .I3(n17781), .O(n836_adj_565[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_10 (.CI(n17743), .I0(n834_adj_574[7]), 
            .I1(n126_c), .CO(n17744));
    SB_LUT4 Error_sub_temp_31__I_0_add_562_9_lut (.I0(Not_Equal_relop1_N_201), 
            .I1(n834_adj_574[6]), .I2(n123_c), .I3(n17742), .O(Switch_out1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_562_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_562_7 (.CI(n17740), .I0(n834_adj_574[4]), 
            .I1(n117_c), .CO(n17741));
    SB_LUT4 add_4257_16_lut (.I0(Not_Equal_relop1_N_201), .I1(n846[14]), 
            .I2(n791_adj_416), .I3(n17725), .O(Switch_out1[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY Error_sub_temp_31__I_0_add_565_3 (.CI(n17781), .I0(n837_adj_572[0]), 
            .I1(n105_c), .CO(n17782));
    SB_CARRY add_4257_16 (.CI(n17725), .I0(n846[14]), .I1(n791_adj_416), 
            .CO(n17726));
    SB_CARRY paramCurrentControlP_15__I_0_add_567_16 (.CI(n17624), .I0(n839[13]), 
            .I1(n761_c), .CO(n763_adj_386));
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_16_lut (.I0(GND_net), .I1(n840[13]), 
            .I2(n765_c), .I3(n17639), .O(n839[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_562_8 (.CI(n17741), .I0(n834_adj_574[5]), 
            .I1(n120_c), .CO(n17742));
    SB_CARRY paramCurrentControlP_15__I_0_add_562_9 (.CI(n17542), .I0(n834[6]), 
            .I1(n102_c), .CO(n17543));
    SB_CARRY Error_sub_temp_31__I_0_add_573_10 (.CI(n17919), .I0(n845_adj_576[7]), 
            .I1(n126_c), .CO(n17920));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_12_lut (.I0(GND_net), .I1(n845_adj_576[9]), 
            .I2(n132_c), .I3(n17921), .O(n844[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4257_15_lut (.I0(Not_Equal_relop1_N_201), .I1(n845_adj_576[14]), 
            .I2(n787_adj_421), .I3(n17724), .O(Switch_out1[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4257_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4257_15 (.CI(n17724), .I0(n845_adj_576[14]), .I1(n787_adj_421), 
            .CO(n17725));
    SB_CARRY paramCurrentControlP_15__I_0_add_568_16 (.CI(n17639), .I0(n840[13]), 
            .I1(n765_c), .CO(n767_adj_382));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_9_lut (.I0(GND_net), .I1(n845_adj_576[6]), 
            .I2(n123_c), .I3(n17918), .O(n844[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_565_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n836_adj_565[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_15_lut (.I0(GND_net), .I1(n840[12]), 
            .I2(n120_c), .I3(n17638), .O(n839[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_9 (.CI(n17918), .I0(n845_adj_576[6]), 
            .I1(n123_c), .CO(n17919));
    SB_CARRY Error_sub_temp_31__I_0_add_565_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17781));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_16_lut (.I0(GND_net), .I1(n836_adj_565[13]), 
            .I2(n146), .I3(n17779), .O(n835_adj_564[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_15 (.CI(n17638), .I0(n840[12]), 
            .I1(n120_c), .CO(n17639));
    SB_CARRY Error_sub_temp_31__I_0_add_564_16 (.CI(n17779), .I0(n836_adj_565[13]), 
            .I1(n146), .CO(n751));
    SB_LUT4 Error_sub_temp_31__I_0_add_564_15_lut (.I0(GND_net), .I1(n836_adj_565[12]), 
            .I2(n141), .I3(n17778), .O(n835_adj_564[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_564_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_564_15 (.CI(n17778), .I0(n836_adj_565[12]), 
            .I1(n141), .CO(n17779));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_8_lut (.I0(GND_net), .I1(n845_adj_576[5]), 
            .I2(n120_c), .I3(n17917), .O(n844[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_14_lut (.I0(GND_net), .I1(n840[11]), 
            .I2(n120_c), .I3(n17637), .O(n839[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_568_14 (.CI(n17637), .I0(n840[11]), 
            .I1(n120_c), .CO(n17638));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_3_lut (.I0(GND_net), .I1(n834[0]), 
            .I2(n102_c), .I3(n17536), .O(n833[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_568_13_lut (.I0(GND_net), .I1(n840[10]), 
            .I2(n120_c), .I3(n17636), .O(n839[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_568_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_8 (.CI(n17917), .I0(n845_adj_576[5]), 
            .I1(n120_c), .CO(n17918));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_7_lut (.I0(GND_net), .I1(n845_adj_576[4]), 
            .I2(n117_c), .I3(n17916), .O(n844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_7 (.CI(n17916), .I0(n845_adj_576[4]), 
            .I1(n117_c), .CO(n17917));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_6_lut (.I0(GND_net), .I1(n845_adj_576[3]), 
            .I2(n114_c), .I3(n17915), .O(n844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_573_6 (.CI(n17915), .I0(n845_adj_576[3]), 
            .I1(n114_c), .CO(n17916));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_5_lut (.I0(GND_net), .I1(n845_adj_576[2]), 
            .I2(n111_c), .I3(n17914), .O(n844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_i61_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[29]), .I2(GND_net), .I3(GND_net), .O(n138_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY Error_sub_temp_31__I_0_add_573_5 (.CI(n17914), .I0(n845_adj_576[2]), 
            .I1(n111_c), .CO(n17915));
    SB_LUT4 add_307_32_lut (.I0(GND_net), .I1(GND_net), .I2(n1[31]), .I3(n15804), 
            .O(\Error_sub_temp[31] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_307_31_lut (.I0(GND_net), .I1(GND_net), .I2(n1[30]), .I3(n15803), 
            .O(\Error_sub_temp[30] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_31 (.CI(n15803), .I0(GND_net), .I1(n1[30]), .CO(n15804));
    SB_LUT4 add_307_30_lut (.I0(GND_net), .I1(GND_net), .I2(n1[29]), .I3(n15802), 
            .O(Error_sub_temp[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Error_sub_temp_31__I_0_add_573_4_lut (.I0(GND_net), .I1(n845_adj_576[1]), 
            .I2(n108_c), .I3(n17913), .O(n844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_30 (.CI(n15802), .I0(GND_net), .I1(n1[29]), .CO(n15803));
    SB_LUT4 add_307_29_lut (.I0(GND_net), .I1(GND_net), .I2(n1[28]), .I3(n15801), 
            .O(Error_sub_temp[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_29 (.CI(n15801), .I0(GND_net), .I1(n1[28]), .CO(n15802));
    SB_LUT4 add_307_28_lut (.I0(GND_net), .I1(GND_net), .I2(n1[27]), .I3(n15800), 
            .O(Error_sub_temp[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_28 (.CI(n15800), .I0(GND_net), .I1(n1[27]), .CO(n15801));
    SB_LUT4 add_307_27_lut (.I0(GND_net), .I1(GND_net), .I2(n1[26]), .I3(n15799), 
            .O(Error_sub_temp[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_27 (.CI(n15799), .I0(GND_net), .I1(n1[26]), .CO(n15800));
    SB_CARRY Error_sub_temp_31__I_0_add_573_4 (.CI(n17913), .I0(n845_adj_576[1]), 
            .I1(n108_c), .CO(n17914));
    SB_LUT4 add_307_26_lut (.I0(GND_net), .I1(GND_net), .I2(n1[25]), .I3(n15798), 
            .O(Error_sub_temp[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_26 (.CI(n15798), .I0(GND_net), .I1(n1[25]), .CO(n15799));
    SB_LUT4 add_307_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[24]), .I3(n15797), 
            .O(Error_sub_temp[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_25 (.CI(n15797), .I0(GND_net), .I1(n1[24]), .CO(n15798));
    SB_LUT4 add_307_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), .I3(n15796), 
            .O(Error_sub_temp[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_24 (.CI(n15796), .I0(GND_net), .I1(n1[23]), .CO(n15797));
    SB_LUT4 add_307_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), .I3(n15795), 
            .O(Error_sub_temp[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_23 (.CI(n15795), .I0(GND_net), .I1(n1[22]), .CO(n15796));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_3_lut (.I0(GND_net), .I1(n845_adj_576[0]), 
            .I2(n105_c), .I3(n17912), .O(n844[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_307_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), .I3(n15794), 
            .O(Error_sub_temp[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_22 (.CI(n15794), .I0(GND_net), .I1(n1[21]), .CO(n15795));
    SB_LUT4 add_307_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), .I3(n15793), 
            .O(Error_sub_temp[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_21 (.CI(n15793), .I0(GND_net), .I1(n1[20]), .CO(n15794));
    SB_LUT4 add_307_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), .I3(n15792), 
            .O(Error_sub_temp[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_20 (.CI(n15792), .I0(GND_net), .I1(n1[19]), .CO(n15793));
    SB_CARRY Error_sub_temp_31__I_0_add_573_3 (.CI(n17912), .I0(n845_adj_576[0]), 
            .I1(n105_c), .CO(n17913));
    SB_LUT4 add_307_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), .I3(n15791), 
            .O(Error_sub_temp[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_19 (.CI(n15791), .I0(GND_net), .I1(n1[18]), .CO(n15792));
    SB_LUT4 add_307_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), .I3(n15790), 
            .O(Error_sub_temp[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_18 (.CI(n15790), .I0(GND_net), .I1(n1[17]), .CO(n15791));
    SB_LUT4 Error_sub_temp_31__I_0_add_573_2_lut (.I0(GND_net), .I1(Proportional_Gain_mul_temp[0]), 
            .I2(n102_c), .I3(GND_net), .O(n844[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_573_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_307_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), .I3(n15789), 
            .O(Error_sub_temp[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_307_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_17 (.CI(n15789), .I0(GND_net), .I1(n1[16]), .CO(n15790));
    SB_CARRY Error_sub_temp_31__I_0_add_573_2 (.CI(GND_net), .I0(Proportional_Gain_mul_temp[0]), 
            .I1(n102_c), .CO(n17912));
    SB_CARRY add_307_16 (.CI(n15788), .I0(GND_net), .I1(n1[15]), .CO(n15789));
    SB_CARRY add_307_15 (.CI(n15787), .I0(GND_net), .I1(n1[14]), .CO(n15788));
    SB_CARRY add_307_14 (.CI(n15786), .I0(GND_net), .I1(n1[13]), .CO(n15787));
    SB_CARRY add_307_13 (.CI(n15785), .I0(GND_net), .I1(n1[12]), .CO(n15786));
    SB_CARRY add_307_12 (.CI(n15784), .I0(GND_net), .I1(n1[11]), .CO(n15785));
    SB_CARRY add_307_11 (.CI(n15783), .I0(GND_net), .I1(n1[10]), .CO(n15784));
    SB_CARRY add_307_10 (.CI(n15782), .I0(GND_net), .I1(n1[9]), .CO(n15783));
    SB_CARRY add_307_9 (.CI(n15781), .I0(GND_net), .I1(n1[8]), .CO(n15782));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_16_lut (.I0(GND_net), .I1(n844[13]), 
            .I2(n146), .I3(n17910), .O(n843[14])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_307_8 (.CI(n15780), .I0(GND_net), .I1(n1[7]), .CO(n15781));
    SB_CARRY add_307_7 (.CI(n15779), .I0(GND_net), .I1(n1[6]), .CO(n15780));
    SB_CARRY add_307_6 (.CI(n15778), .I0(GND_net), .I1(n1[5]), .CO(n15779));
    SB_CARRY add_307_5 (.CI(n15777), .I0(GND_net), .I1(n1[4]), .CO(n15778));
    SB_CARRY add_307_4 (.CI(n15776), .I0(GND_net), .I1(n1[3]), .CO(n15777));
    SB_CARRY add_307_3 (.CI(n15775), .I0(GND_net), .I1(n31), .CO(n15776));
    SB_CARRY add_307_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n15775));
    SB_CARRY Error_sub_temp_31__I_0_add_572_16 (.CI(n17910), .I0(n844[13]), 
            .I1(n146), .CO(n783));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_15_lut (.I0(GND_net), .I1(n844[12]), 
            .I2(n141), .I3(n17909), .O(n843[13])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_add_566_16_lut (.I0(GND_net), .I1(n838[13]), 
            .I2(n757_c), .I3(n17609), .O(n837[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_566_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_15 (.CI(n17909), .I0(n844[12]), 
            .I1(n141), .CO(n17910));
    SB_LUT4 paramCurrentControlP_15__I_0_i49_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[23]), .I2(GND_net), .I3(GND_net), .O(n120_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i49_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i41_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[19]), .I2(GND_net), .I3(GND_net), .O(n108_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i41_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i47_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[22]), .I2(GND_net), .I3(GND_net), .O(n117_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i47_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i39_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[18]), .I2(GND_net), .I3(GND_net), .O(n105_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i39_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i513_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[21]), .I2(GND_net), .I3(GND_net), .O(n757_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i513_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i45_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[21]), .I2(GND_net), .I3(GND_net), .O(n114_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i45_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i35_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[16]), .I2(GND_net), .I3(GND_net), .O(Proportional_Gain_mul_temp[0]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i35_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Error_sub_temp_31__I_0_add_572_14_lut (.I0(GND_net), .I1(n844[11]), 
            .I2(n138_c), .I3(n17908), .O(n843[12])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_14 (.CI(n17908), .I0(n844[11]), 
            .I1(n138_c), .CO(n17909));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_13_lut (.I0(GND_net), .I1(n844[10]), 
            .I2(n135_c), .I3(n17907), .O(n843[11])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_13 (.CI(n17907), .I0(n844[10]), 
            .I1(n135_c), .CO(n17908));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_12_lut (.I0(GND_net), .I1(n844[9]), 
            .I2(n132_c), .I3(n17906), .O(n843[10])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_12 (.CI(n17906), .I0(n844[9]), 
            .I1(n132_c), .CO(n17907));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_11_lut (.I0(GND_net), .I1(n844[8]), 
            .I2(n129_c), .I3(n17905), .O(n843[9])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF currentControlITerm_i4 (.Q(currentControlITerm[4]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14323));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_CARRY Error_sub_temp_31__I_0_add_572_11 (.CI(n17905), .I0(n844[8]), 
            .I1(n129_c), .CO(n17906));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_10_lut (.I0(GND_net), .I1(n844[7]), 
            .I2(n126_c), .I3(n17904), .O(n843[8])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_10 (.CI(n17904), .I0(n844[7]), 
            .I1(n126_c), .CO(n17905));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_9_lut (.I0(GND_net), .I1(n844[6]), 
            .I2(n123_c), .I3(n17903), .O(n843[7])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF currentControlITerm_i2 (.Q(currentControlITerm[2]), .C(pin3_clk_16mhz_N_keep), 
           .D(n14321));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(127[10] 137[8])
    SB_CARRY Error_sub_temp_31__I_0_add_572_9 (.CI(n17903), .I0(n844[6]), 
            .I1(n123_c), .CO(n17904));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_8_lut (.I0(GND_net), .I1(n844[5]), 
            .I2(n120_c), .I3(n17902), .O(n843[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_8 (.CI(n17902), .I0(n844[5]), 
            .I1(n120_c), .CO(n17903));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_7_lut (.I0(GND_net), .I1(n844[4]), 
            .I2(n117_c), .I3(n17901), .O(n843[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Error_sub_temp_31__I_0_add_572_7 (.CI(n17901), .I0(n844[4]), 
            .I1(n117_c), .CO(n17902));
    SB_CARRY paramCurrentControlP_15__I_0_add_568_13 (.CI(n17636), .I0(n840[10]), 
            .I1(n120_c), .CO(n17637));
    SB_LUT4 Error_sub_temp_31__I_0_add_572_4_lut (.I0(GND_net), .I1(n844[1]), 
            .I2(n108_c), .I3(n17898), .O(n843[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Error_sub_temp_31__I_0_add_572_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 paramCurrentControlP_15__I_0_i528_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[26]), .I2(GND_net), .I3(GND_net), .O(n777_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i528_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i43_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[20]), .I2(GND_net), .I3(GND_net), .O(n111_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i43_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_i55_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[26]), .I2(GND_net), .I3(GND_net), .O(n129_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_130 (.I0(\Add_add_temp[5] ), .I1(\Add_add_temp[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n20712));
    defparam i1_2_lut_adj_130.LUT_INIT = 16'h8888;
    SB_LUT4 paramCurrentControlP_15__I_0_add_569_16_lut (.I0(GND_net), .I1(n841[11]), 
            .I2(n769_c), .I3(n17654), .O(n840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_569_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_3 (.CI(n17536), .I0(n834[0]), 
            .I1(n102_c), .CO(n17537));
    SB_LUT4 paramCurrentControlP_15__I_0_add_562_2_lut (.I0(GND_net), .I1(n105_c), 
            .I2(n102_c), .I3(GND_net), .O(n833[0])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_562_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_562_2 (.CI(GND_net), .I0(n105_c), 
            .I1(n102_c), .CO(n17536));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_16_lut (.I0(GND_net), .I1(n833[13]), 
            .I2(n737_c), .I3(n17534), .O(n832[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_16 (.CI(n17534), .I0(n833[13]), 
            .I1(n737_c), .CO(n739));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_15_lut (.I0(GND_net), .I1(n833[12]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17533), .O(Proportional_Gain_mul_temp[14])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_15 (.CI(n17533), .I0(n833[12]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17534));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_14_lut (.I0(GND_net), .I1(n833[11]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17532), .O(Proportional_Gain_mul_temp[13])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_14 (.CI(n17532), .I0(n833[11]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17533));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_13_lut (.I0(GND_net), .I1(n833[10]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17531), .O(Proportional_Gain_mul_temp[12])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_13 (.CI(n17531), .I0(n833[10]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17532));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_12_lut (.I0(GND_net), .I1(n833[9]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17530), .O(Proportional_Gain_mul_temp[11])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_12 (.CI(n17530), .I0(n833[9]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17531));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_11_lut (.I0(GND_net), .I1(n833[8]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17529), .O(Proportional_Gain_mul_temp[10])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_11 (.CI(n17529), .I0(n833[8]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17530));
    SB_LUT4 paramCurrentControlP_15__I_0_add_563_3_lut (.I0(GND_net), .I1(n835[0]), 
            .I2(n105_c), .I3(n17551), .O(n834[1])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_131 (.I0(\Add_add_temp[7] ), .I1(\Add_add_temp[8] ), 
            .I2(\Add_add_temp[6] ), .I3(n20712), .O(n19777));
    defparam i1_4_lut_adj_131.LUT_INIT = 16'h8000;
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_10_lut (.I0(GND_net), .I1(n833[7]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17528), .O(Proportional_Gain_mul_temp[9])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_10 (.CI(n17528), .I0(n833[7]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17529));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_9_lut (.I0(GND_net), .I1(n833[6]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17527), .O(Proportional_Gain_mul_temp[8])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY paramCurrentControlP_15__I_0_add_561_9 (.CI(n17527), .I0(n833[6]), 
            .I1(Proportional_Gain_mul_temp[0]), .CO(n17528));
    SB_LUT4 paramCurrentControlP_15__I_0_add_561_8_lut (.I0(GND_net), .I1(n833[5]), 
            .I2(Proportional_Gain_mul_temp[0]), .I3(n17526), .O(Proportional_Gain_mul_temp[7])) /* synthesis syn_instantiated=1 */ ;
    defparam paramCurrentControlP_15__I_0_add_561_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_132 (.I0(\Add_add_temp[11] ), .I1(n19777), .I2(\Add_add_temp[10] ), 
            .I3(\Add_add_temp[9] ), .O(n20700));
    defparam i1_4_lut_adj_132.LUT_INIT = 16'hfaea;
    SB_LUT4 i13268_4_lut (.I0(\Add_add_temp[12] ), .I1(\Add_add_temp[14] ), 
            .I2(\Add_add_temp[13] ), .I3(n20700), .O(n15205));
    defparam i13268_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut_adj_133 (.I0(\Add_add_temp[17] ), .I1(n15205), .I2(\Add_add_temp[16] ), 
            .I3(\Add_add_temp[15] ), .O(n20670));
    defparam i1_4_lut_adj_133.LUT_INIT = 16'hfaea;
    SB_LUT4 i1_4_lut_adj_134 (.I0(\Add_add_temp[19] ), .I1(\Add_add_temp[20] ), 
            .I2(\Add_add_temp[18] ), .I3(n20670), .O(n19746));
    defparam i1_4_lut_adj_134.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_135 (.I0(n19269), .I1(n789_c), .I2(n19273), .I3(n142), 
            .O(n845[14]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_4_lut_adj_135.LUT_INIT = 16'hc966;
    SB_LUT4 i1_4_lut_adj_136 (.I0(\Add_add_temp[23] ), .I1(n19746), .I2(\Add_add_temp[22] ), 
            .I3(\Add_add_temp[21] ), .O(n20656));
    defparam i1_4_lut_adj_136.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_137 (.I0(\Add_add_temp[26] ), .I1(n20656), .I2(\Add_add_temp[25] ), 
            .I3(\Add_add_temp[24] ), .O(n20648));
    defparam i1_4_lut_adj_137.LUT_INIT = 16'hfaea;
    SB_LUT4 i1_4_lut_adj_138 (.I0(\Add_add_temp[29] ), .I1(n20648), .I2(\Add_add_temp[28] ), 
            .I3(\Add_add_temp[27] ), .O(n20634));
    defparam i1_4_lut_adj_138.LUT_INIT = 16'hfaea;
    SB_LUT4 i13327_4_lut (.I0(\Add_add_temp[30] ), .I1(\Add_add_temp[32] ), 
            .I2(\Add_add_temp[31] ), .I3(n20634), .O(n15264));
    defparam i13327_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut_adj_139 (.I0(\Add_add_temp[34] ), .I1(Saturate_out1[31]), 
            .I2(\Add_add_temp[33] ), .I3(n15264), .O(Saturate_out1_31__N_267));
    defparam i1_4_lut_adj_139.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_140 (.I0(\Add_add_temp[7] ), .I1(\Add_add_temp[8] ), 
            .I2(\Add_add_temp[6] ), .I3(\Add_add_temp[5] ), .O(n19723));
    defparam i1_4_lut_adj_140.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_141 (.I0(\Add_add_temp[11] ), .I1(n19723), .I2(\Add_add_temp[10] ), 
            .I3(\Add_add_temp[9] ), .O(n20708));
    defparam i1_4_lut_adj_141.LUT_INIT = 16'ha8a0;
    SB_LUT4 i729_4_lut (.I0(\Add_add_temp[12] ), .I1(\Add_add_temp[14] ), 
            .I2(\Add_add_temp[13] ), .I3(n20708), .O(n22_adj_519));
    defparam i729_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_142 (.I0(\Add_add_temp[17] ), .I1(n22_adj_519), 
            .I2(\Add_add_temp[16] ), .I3(\Add_add_temp[15] ), .O(n20688));
    defparam i1_4_lut_adj_142.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_143 (.I0(\Add_add_temp[19] ), .I1(\Add_add_temp[20] ), 
            .I2(\Add_add_temp[18] ), .I3(n20688), .O(n19842));
    defparam i1_4_lut_adj_143.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_144 (.I0(\Add_add_temp[23] ), .I1(n19842), .I2(\Add_add_temp[22] ), 
            .I3(\Add_add_temp[21] ), .O(n20666));
    defparam i1_4_lut_adj_144.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_145 (.I0(\Add_add_temp[26] ), .I1(n20666), .I2(\Add_add_temp[25] ), 
            .I3(\Add_add_temp[24] ), .O(n20658));
    defparam i1_4_lut_adj_145.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_146 (.I0(\Add_add_temp[29] ), .I1(n20658), .I2(\Add_add_temp[28] ), 
            .I3(\Add_add_temp[27] ), .O(n20644));
    defparam i1_4_lut_adj_146.LUT_INIT = 16'ha8a0;
    SB_LUT4 i747_4_lut (.I0(\Add_add_temp[30] ), .I1(\Add_add_temp[32] ), 
            .I2(\Add_add_temp[31] ), .I3(n20644), .O(n58));
    defparam i747_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_147 (.I0(\Add_add_temp[34] ), .I1(Saturate_out1[31]), 
            .I2(\Add_add_temp[33] ), .I3(n58), .O(Saturate_out1_31__N_266));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(121[27:75])
    defparam i1_4_lut_adj_147.LUT_INIT = 16'h2000;
    SB_LUT4 paramCurrentControlP_15__I_0_i57_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[27]), .I2(GND_net), .I3(GND_net), .O(n132_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_76_inv_0_i4_1_lut (.I0(\dCurrent[3] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i5_1_lut (.I0(\dCurrent[4] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i6_1_lut (.I0(\dCurrent[5] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i7_1_lut (.I0(\dCurrent[6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i8_1_lut (.I0(\dCurrent[7] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i9_1_lut (.I0(\dCurrent[8] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i10_1_lut (.I0(\dCurrent[9] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[9]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i11_1_lut (.I0(\dCurrent[10] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[10]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i12_1_lut (.I0(\dCurrent[11] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[11]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i13_1_lut (.I0(\dCurrent[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[12]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i14_1_lut (.I0(\dCurrent[13] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[13]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i15_1_lut (.I0(\dCurrent[14] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[14]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i16_1_lut (.I0(\dCurrent[15] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[15]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i17_1_lut (.I0(\dCurrent[16] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[16]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i18_1_lut (.I0(\dCurrent[17] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[17]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i19_1_lut (.I0(\dCurrent[18] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[18]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i20_1_lut (.I0(\dCurrent[19] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[19]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i21_1_lut (.I0(\dCurrent[20] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[20]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i22_1_lut (.I0(\dCurrent[21] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[21]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i23_1_lut (.I0(\dCurrent[22] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[22]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 paramCurrentControlP_15__I_0_i53_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[25]), .I2(GND_net), .I3(GND_net), .O(n126_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_76_inv_0_i24_1_lut (.I0(\dCurrent[23] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[23]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i25_1_lut (.I0(\dCurrent[24] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[24]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i26_1_lut (.I0(\dCurrent[25] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[25]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i27_1_lut (.I0(\dCurrent[26] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[26]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i28_1_lut (.I0(\dCurrent[27] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[27]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i29_1_lut (.I0(\dCurrent[28] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[28]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i30_1_lut (.I0(\dCurrent[29] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[29]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i31_1_lut (.I0(\dCurrent[30] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[30]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_76_inv_0_i32_1_lut (.I0(\dCurrent[31] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[31]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(73[27:60])
    defparam sub_76_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6570_2_lut (.I0(n833_adj_575[13]), .I1(\Error_sub_temp[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n832_adj_577[14]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(92[30:64])
    defparam i6570_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 paramCurrentControlP_15__I_0_i498_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[16]), .I2(GND_net), .I3(GND_net), .O(n737_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i498_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i501_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[17]), .I2(GND_net), .I3(GND_net), .O(n741_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i501_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i504_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[18]), .I2(GND_net), .I3(GND_net), .O(n745_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i504_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i507_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[19]), .I2(GND_net), .I3(GND_net), .O(n749_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i507_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i510_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[20]), .I2(GND_net), .I3(GND_net), .O(n753_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i510_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i516_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[22]), .I2(GND_net), .I3(GND_net), .O(n761_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i516_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i519_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[23]), .I2(GND_net), .I3(GND_net), .O(n765_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i519_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_3_lut (.I0(n138_c), .I1(n142), .I2(n12), .I3(n12), 
            .O(n19273));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_4_lut_3_lut.LUT_INIT = 16'heeaa;
    SB_LUT4 paramCurrentControlP_15__I_0_i525_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[25]), .I2(GND_net), .I3(GND_net), .O(n773_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i525_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 paramCurrentControlP_15__I_0_i531_2_lut (.I0(\Product_mul_temp[26] ), 
            .I1(Error_sub_temp[27]), .I2(GND_net), .I3(GND_net), .O(n781_c));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam paramCurrentControlP_15__I_0_i531_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_4_lut (.I0(n142), .I1(\Product_mul_temp[26] ), 
            .I2(Error_sub_temp[29]), .I3(n4), .O(n12));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_2_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Product_mul_temp[26] ), .I1(Error_sub_temp[29]), 
            .I2(n142), .I3(n4), .O(n845[3]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h80f8;
    SB_LUT4 i2_3_lut_4_lut (.I0(n4), .I1(\Product_mul_temp[26] ), .I2(Error_sub_temp[29]), 
            .I3(n142), .O(n845[2]));   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(78[39:81])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h956a;
    Saturate_Output_U0 u_Saturate_Output (.\preSatVoltage[15] (preSatVoltage[15]), 
            .Out_31__N_333(Out_31__N_333), .\Product_mul_temp[26] (\Product_mul_temp[26] ), 
            .Out_31__N_332(Out_31__N_332), .n342(n342), .\dVoltage[6] (\dVoltage[6] ), 
            .GND_net(GND_net), .Look_Up_Table_out1_1({Look_Up_Table_out1_1}), 
            .n342_adj_1(n342_adj_10), .\preSatVoltage[11] (preSatVoltage[11]), 
            .n114(n114), .\preSatVoltage[17] (preSatVoltage[17]), .\preSatVoltage[16] (preSatVoltage[16]), 
            .\preSatVoltage[19] (\preSatVoltage[19] ), .\preSatVoltage[20] (preSatVoltage[20]), 
            .\preSatVoltage[18] (preSatVoltage[18]), .n408(n408), .\preSatVoltage[9] (preSatVoltage[9]), 
            .n14(n14), .n20198(n20198), .\preSatVoltage[10] (\preSatVoltage[10] ), 
            .\preSatVoltage[21] (preSatVoltage[21]), .n604(n604), .\preSatVoltage[12] (\preSatVoltage[12] ), 
            .\preSatVoltage[13] (preSatVoltage[13]), .\preSatVoltage[22] (preSatVoltage[22]), 
            .n685(n685), .n685_adj_2(n685_adj_11), .\dVoltage[13] (\dVoltage[13] ), 
            .\preSatVoltage[14] (preSatVoltage[14]), .n417(n417), .n123(n123), 
            .\preSatVoltage[25] (preSatVoltage[25]), .\preSatVoltage[24] (preSatVoltage[24]), 
            .\preSatVoltage[23] (\preSatVoltage[23] ), .\preSatVoltage[28] (preSatVoltage[28]), 
            .\preSatVoltage[27] (preSatVoltage[27]), .\preSatVoltage[26] (preSatVoltage[26]), 
            .n613(n613), .n429(n429), .\preSatVoltage[29] (preSatVoltage[29]), 
            .\Voltage_1[31] (Voltage_1[31]), .\preSatVoltage[30] (preSatVoltage[30]), 
            .n135(n135), .n625(n625), .n587(n587), .n587_adj_3(n587_adj_12), 
            .\dVoltage[11] (\dVoltage[11] ), .n399(n399), .n426(n426), 
            .n414(n414), .n432(n432), .n393(n393), .n405(n405), .n402(n402), 
            .n396(n396), .n420(n420), .n423(n423), .\dVoltage[8] (\dVoltage[8] ), 
            .n44(n44), .n489(n489), .n8(n8), .\dVoltage[9] (\dVoltage[9] ), 
            .n489_adj_4(n489_adj_13), .n20(n20), .n126(n126), .n616(n616), 
            .n391(n391), .\dVoltage[7] (\dVoltage[7] ), .n391_adj_5(n391_adj_14), 
            .n19576(n19576), .n129(n129), .n619(n619), .n11(n11), .n35(n35), 
            .n19352(n19352), .n26(n26), .\Product3_mul_temp[2] (\Product3_mul_temp[2] ), 
            .n120(n120), .n111(n111), .n102(n102), .n99(n99), .n108(n108), 
            .n138(n138), .n132(n132), .n105(n105), .\dVoltage[2] (\dVoltage[2] ), 
            .n610(n610), .n595(n595), .n23(n23), .n622(n622), .n41(n41), 
            .n601(n601), .n592(n592), .n598(n598), .n589(n589), .n628(n628), 
            .n32(n32), .\dVoltage[12] (\dVoltage[12] ), .\dVoltage[10] (\dVoltage[10] ), 
            .n538(n538), .n29(n29), .n17(n17), .n71(n71), .n83(n83), 
            .n59(n59), .n50(n50), .n92(n92), .n68(n68), .n62(n62), 
            .n53(n53), .n65(n65), .n38(n38), .n56(n56), .n80(n80), 
            .n244(n244), .n233(n233), .n14_adj_6(n14_c), .n200(n200), 
            .n203(n203), .n86(n86), .n77(n77), .n197(n197), .n239(n239), 
            .n206(n206), .n86_adj_7(n86_adj_15), .n215(n215), .n89(n89), 
            .n74(n74), .n227(n227), .n233_adj_8(n233_adj_16), .n224(n224), 
            .n221(n221), .n209(n209), .n236(n236), .n230(n230), .n244_adj_9(n244_adj_17), 
            .n212(n212), .n218(n218), .n279(n279), .n270(n270), .n267(n267), 
            .n255(n255), .n285(n285), .n264(n264), .n258(n258), .n249(n249), 
            .n246(n246), .n273(n273), .\dVoltage[14] (\dVoltage[14] ), 
            .n282(n282), .n261(n261), .n19681(n19681), .n288(n288), 
            .n276(n276), .n252(n252), .\dVoltage[5] (\dVoltage[5] ), .n789(n789), 
            .n785(n785), .n765(n765), .n753(n753), .n741(n741), .n757(n757), 
            .n745(n745), .n761(n761), .n195(n195), .n737(n737), .\dVoltage[3] (\dVoltage[3] ), 
            .n749(n749), .n781(n781), .n777(n777), .n773(n773), .n769(n769), 
            .n19684(n19684), .\dVoltage[15] (\dVoltage[15] ), .n435(n435), 
            .n141(n141_adj_18), .n631(n631), .n117(n117), .n411(n411), 
            .n607(n607)) /* synthesis syn_module_defined=1 */ ;   // ../../hdlcoderFocCurrentFixptHdl/D_Current_Control.v(148[19] 150[39])
    VCC i1 (.Y(VCC_net));
    
endmodule
//
// Verilog Description of module Saturate_Output_U0
//

module Saturate_Output_U0 (\preSatVoltage[15] , Out_31__N_333, \Product_mul_temp[26] , 
            Out_31__N_332, n342, \dVoltage[6] , GND_net, Look_Up_Table_out1_1, 
            n342_adj_1, \preSatVoltage[11] , n114, \preSatVoltage[17] , 
            \preSatVoltage[16] , \preSatVoltage[19] , \preSatVoltage[20] , 
            \preSatVoltage[18] , n408, \preSatVoltage[9] , n14, n20198, 
            \preSatVoltage[10] , \preSatVoltage[21] , n604, \preSatVoltage[12] , 
            \preSatVoltage[13] , \preSatVoltage[22] , n685, n685_adj_2, 
            \dVoltage[13] , \preSatVoltage[14] , n417, n123, \preSatVoltage[25] , 
            \preSatVoltage[24] , \preSatVoltage[23] , \preSatVoltage[28] , 
            \preSatVoltage[27] , \preSatVoltage[26] , n613, n429, \preSatVoltage[29] , 
            \Voltage_1[31] , \preSatVoltage[30] , n135, n625, n587, 
            n587_adj_3, \dVoltage[11] , n399, n426, n414, n432, 
            n393, n405, n402, n396, n420, n423, \dVoltage[8] , 
            n44, n489, n8, \dVoltage[9] , n489_adj_4, n20, n126, 
            n616, n391, \dVoltage[7] , n391_adj_5, n19576, n129, 
            n619, n11, n35, n19352, n26, \Product3_mul_temp[2] , 
            n120, n111, n102, n99, n108, n138, n132, n105, \dVoltage[2] , 
            n610, n595, n23, n622, n41, n601, n592, n598, n589, 
            n628, n32, \dVoltage[12] , \dVoltage[10] , n538, n29, 
            n17, n71, n83, n59, n50, n92, n68, n62, n53, n65, 
            n38, n56, n80, n244, n233, n14_adj_6, n200, n203, 
            n86, n77, n197, n239, n206, n86_adj_7, n215, n89, 
            n74, n227, n233_adj_8, n224, n221, n209, n236, n230, 
            n244_adj_9, n212, n218, n279, n270, n267, n255, n285, 
            n264, n258, n249, n246, n273, \dVoltage[14] , n282, 
            n261, n19681, n288, n276, n252, \dVoltage[5] , n789, 
            n785, n765, n753, n741, n757, n745, n761, n195, 
            n737, \dVoltage[3] , n749, n781, n777, n773, n769, 
            n19684, \dVoltage[15] , n435, n141, n631, n117, n411, 
            n607) /* synthesis syn_module_defined=1 */ ;
    input \preSatVoltage[15] ;
    output Out_31__N_333;
    input \Product_mul_temp[26] ;
    output Out_31__N_332;
    output n342;
    output \dVoltage[6] ;
    input GND_net;
    input [15:0]Look_Up_Table_out1_1;
    output n342_adj_1;
    input \preSatVoltage[11] ;
    output n114;
    input \preSatVoltage[17] ;
    input \preSatVoltage[16] ;
    input \preSatVoltage[19] ;
    input \preSatVoltage[20] ;
    input \preSatVoltage[18] ;
    output n408;
    input \preSatVoltage[9] ;
    output n14;
    input n20198;
    input \preSatVoltage[10] ;
    input \preSatVoltage[21] ;
    output n604;
    input \preSatVoltage[12] ;
    input \preSatVoltage[13] ;
    input \preSatVoltage[22] ;
    output n685;
    output n685_adj_2;
    output \dVoltage[13] ;
    input \preSatVoltage[14] ;
    output n417;
    output n123;
    input \preSatVoltage[25] ;
    input \preSatVoltage[24] ;
    input \preSatVoltage[23] ;
    input \preSatVoltage[28] ;
    input \preSatVoltage[27] ;
    input \preSatVoltage[26] ;
    output n613;
    output n429;
    input \preSatVoltage[29] ;
    input \Voltage_1[31] ;
    input \preSatVoltage[30] ;
    output n135;
    output n625;
    output n587;
    output n587_adj_3;
    output \dVoltage[11] ;
    output n399;
    output n426;
    output n414;
    output n432;
    output n393;
    output n405;
    output n402;
    output n396;
    output n420;
    output n423;
    output \dVoltage[8] ;
    output n44;
    output n489;
    output n8;
    output \dVoltage[9] ;
    output n489_adj_4;
    output n20;
    output n126;
    output n616;
    output n391;
    output \dVoltage[7] ;
    output n391_adj_5;
    output n19576;
    output n129;
    output n619;
    output n11;
    output n35;
    output n19352;
    output n26;
    output \Product3_mul_temp[2] ;
    output n120;
    output n111;
    output n102;
    output n99;
    output n108;
    output n138;
    output n132;
    output n105;
    output \dVoltage[2] ;
    output n610;
    output n595;
    output n23;
    output n622;
    output n41;
    output n601;
    output n592;
    output n598;
    output n589;
    output n628;
    output n32;
    output \dVoltage[12] ;
    output \dVoltage[10] ;
    output n538;
    output n29;
    output n17;
    output n71;
    output n83;
    output n59;
    output n50;
    output n92;
    output n68;
    output n62;
    output n53;
    output n65;
    output n38;
    output n56;
    output n80;
    output n244;
    output n233;
    output n14_adj_6;
    output n200;
    output n203;
    output n86;
    output n77;
    output n197;
    output n239;
    output n206;
    output n86_adj_7;
    output n215;
    output n89;
    output n74;
    output n227;
    output n233_adj_8;
    output n224;
    output n221;
    output n209;
    output n236;
    output n230;
    output n244_adj_9;
    output n212;
    output n218;
    output n279;
    output n270;
    output n267;
    output n255;
    output n285;
    output n264;
    output n258;
    output n249;
    output n246;
    output n273;
    output \dVoltage[14] ;
    output n282;
    output n261;
    output n19681;
    output n288;
    output n276;
    output n252;
    output \dVoltage[5] ;
    output n789;
    output n785;
    output n765;
    output n753;
    output n741;
    output n757;
    output n745;
    output n761;
    output n195;
    output n737;
    output \dVoltage[3] ;
    output n749;
    output n781;
    output n777;
    output n773;
    output n769;
    output n19684;
    output \dVoltage[15] ;
    output n435;
    output n141;
    output n631;
    output n117;
    output n411;
    output n607;
    
    
    wire n15171, n15188, n19688, n22, n19455, n19690, n20112, 
        n20098, n19926, n19932, n19424, n14851, n19904, n19747;
    
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\preSatVoltage[15] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n342));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h00d0;
    SB_LUT4 i13165_2_lut_3_lut (.I0(\preSatVoltage[15] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[6] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13165_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_7 (.I0(\preSatVoltage[15] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n342_adj_1));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_7.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_8 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[5]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n114));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_8.LUT_INIT = 16'h4440;
    SB_LUT4 i13251_4_lut (.I0(\preSatVoltage[15] ), .I1(\preSatVoltage[17] ), 
            .I2(\preSatVoltage[16] ), .I3(n15171), .O(n15188));
    defparam i13251_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_4_lut (.I0(\preSatVoltage[19] ), .I1(\preSatVoltage[20] ), 
            .I2(\preSatVoltage[18] ), .I3(n15188), .O(n19688));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_9 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[5]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n408));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_9.LUT_INIT = 16'h4440;
    SB_LUT4 i3_4_lut (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), .I2(Out_31__N_333), 
            .I3(Look_Up_Table_out1_1[4]), .O(n14));
    defparam i3_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1202_3_lut (.I0(n20198), .I1(\preSatVoltage[10] ), .I2(\preSatVoltage[9] ), 
            .I3(GND_net), .O(n22));
    defparam i1202_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_10 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[5]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n604));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_10.LUT_INIT = 16'h4440;
    SB_LUT4 i1_4_lut_adj_11 (.I0(\preSatVoltage[12] ), .I1(\preSatVoltage[13] ), 
            .I2(n22), .I3(\preSatVoltage[11] ), .O(n19455));
    defparam i1_4_lut_adj_11.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.I0(\preSatVoltage[22] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n685));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_12.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.I0(\preSatVoltage[22] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n685_adj_2));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_13.LUT_INIT = 16'h00d0;
    SB_LUT4 i13172_2_lut_3_lut (.I0(\preSatVoltage[22] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[13] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13172_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_4_lut_adj_14 (.I0(\preSatVoltage[15] ), .I1(\preSatVoltage[16] ), 
            .I2(n19455), .I3(\preSatVoltage[14] ), .O(n19690));
    defparam i1_4_lut_adj_14.LUT_INIT = 16'h8880;
    SB_LUT4 i1_4_lut_adj_15 (.I0(\preSatVoltage[19] ), .I1(\preSatVoltage[18] ), 
            .I2(n19690), .I3(\preSatVoltage[17] ), .O(n20112));
    defparam i1_4_lut_adj_15.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[8]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n417));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_16.LUT_INIT = 16'h4440;
    SB_LUT4 i1_4_lut_adj_17 (.I0(\preSatVoltage[22] ), .I1(n20112), .I2(\preSatVoltage[21] ), 
            .I3(\preSatVoltage[20] ), .O(n20098));
    defparam i1_4_lut_adj_17.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_18 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[8]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n123));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_18.LUT_INIT = 16'h4440;
    SB_LUT4 i1_4_lut_adj_19 (.I0(\preSatVoltage[25] ), .I1(\preSatVoltage[24] ), 
            .I2(n20098), .I3(\preSatVoltage[23] ), .O(n19926));
    defparam i1_4_lut_adj_19.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_20 (.I0(\preSatVoltage[28] ), .I1(\preSatVoltage[27] ), 
            .I2(\preSatVoltage[26] ), .I3(n19926), .O(n19932));
    defparam i1_4_lut_adj_20.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_21 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[8]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n613));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_21.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_22 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[12]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n429));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_22.LUT_INIT = 16'h4440;
    SB_LUT4 i12820_4_lut (.I0(\preSatVoltage[29] ), .I1(\Voltage_1[31] ), 
            .I2(\preSatVoltage[30] ), .I3(n19932), .O(Out_31__N_332));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[37:72])
    defparam i12820_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[12]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n135));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_23.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_24 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[12]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n625));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_24.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_25 (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n587));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_25.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_26 (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n587_adj_3));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_26.LUT_INIT = 16'h00d0;
    SB_LUT4 i13170_2_lut_3_lut (.I0(\preSatVoltage[20] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[11] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13170_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_4_lut_adj_27 (.I0(\preSatVoltage[22] ), .I1(\preSatVoltage[23] ), 
            .I2(n19688), .I3(\preSatVoltage[21] ), .O(n19424));
    defparam i1_4_lut_adj_27.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n399));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_28.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_29 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n426));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_29.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_30 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), .O(n414));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_30.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_31 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n432));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_31.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_32 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n393));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_32.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_33 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n405));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_33.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n402));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_34.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_35 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n396));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_35.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), .O(n420));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_36.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_37 (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), .O(n423));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_37.LUT_INIT = 16'h00e0;
    SB_LUT4 i13167_2_lut_3_lut (.I0(\preSatVoltage[17] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[8] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13167_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i3_4_lut_adj_38 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[14]), .O(n44));
    defparam i3_4_lut_adj_38.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_39 (.I0(\preSatVoltage[18] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n489));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_39.LUT_INIT = 16'h00d0;
    SB_LUT4 i3_4_lut_adj_40 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[2]), .O(n8));
    defparam i3_4_lut_adj_40.LUT_INIT = 16'h0400;
    SB_LUT4 i13168_2_lut_3_lut (.I0(\preSatVoltage[18] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[9] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13168_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_41 (.I0(\preSatVoltage[18] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n489_adj_4));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_41.LUT_INIT = 16'h00d0;
    SB_LUT4 i3_4_lut_adj_42 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[6]), .O(n20));
    defparam i3_4_lut_adj_42.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[9]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n126));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_43.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[9]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n616));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_44.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_45 (.I0(\preSatVoltage[16] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n391));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_45.LUT_INIT = 16'h00d0;
    SB_LUT4 i13166_2_lut_3_lut (.I0(\preSatVoltage[16] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[7] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13166_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.I0(\preSatVoltage[16] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n391_adj_5));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_46.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_4_lut_adj_47 (.I0(Out_31__N_332), .I1(Out_31__N_333), .I2(\preSatVoltage[9] ), 
            .I3(Look_Up_Table_out1_1[1]), .O(n19576));
    defparam i1_4_lut_adj_47.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_48 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[10]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n129));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_48.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_49 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[10]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n619));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_49.LUT_INIT = 16'h4440;
    SB_LUT4 i3_4_lut_adj_50 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[3]), .O(n11));
    defparam i3_4_lut_adj_50.LUT_INIT = 16'h0400;
    SB_LUT4 i3_4_lut_adj_51 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[11]), .O(n35));
    defparam i3_4_lut_adj_51.LUT_INIT = 16'h0400;
    SB_LUT4 i12876_rep_4_3_lut (.I0(\preSatVoltage[9] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(n19352));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i12876_rep_4_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i3_4_lut_adj_52 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[8]), .O(n26));
    defparam i3_4_lut_adj_52.LUT_INIT = 16'h0400;
    SB_LUT4 i13232_4_lut (.I0(\preSatVoltage[12] ), .I1(\preSatVoltage[14] ), 
            .I2(\preSatVoltage[13] ), .I3(n14851), .O(n15171));
    defparam i13232_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i12921_2_lut (.I0(\preSatVoltage[10] ), .I1(\preSatVoltage[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n14851));
    defparam i12921_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\preSatVoltage[28] ), .I1(\preSatVoltage[27] ), 
            .I2(\preSatVoltage[26] ), .I3(GND_net), .O(n19904));
    defparam i1_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_53 (.I0(\preSatVoltage[25] ), .I1(\preSatVoltage[29] ), 
            .I2(\preSatVoltage[24] ), .I3(n19424), .O(n19747));
    defparam i1_4_lut_adj_53.LUT_INIT = 16'h8000;
    SB_LUT4 i1212_rep_6_4_lut (.I0(n19747), .I1(\Voltage_1[31] ), .I2(\preSatVoltage[30] ), 
            .I3(n19904), .O(Out_31__N_333));
    defparam i1212_rep_6_4_lut.LUT_INIT = 16'h4ccc;
    SB_LUT4 i3_4_lut_adj_54 (.I0(Out_31__N_332), .I1(Out_31__N_333), .I2(\preSatVoltage[9] ), 
            .I3(\Product_mul_temp[26] ), .O(\Product3_mul_temp[2] ));
    defparam i3_4_lut_adj_54.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_55 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), .O(n120));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_55.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_56 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n111));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_56.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_57 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n102));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_57.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n99));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_58.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n108));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_59.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n138));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_60.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n132));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_61.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_62 (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n105));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_62.LUT_INIT = 16'h00e0;
    SB_LUT4 i13161_2_lut_3_lut (.I0(\preSatVoltage[11] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[2] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13161_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_63 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[7]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n610));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_63.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_64 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n595));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_64.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_65 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[7]), .O(n23));
    defparam i3_4_lut_adj_65.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_66 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n622));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_66.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_67 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[13]), .O(n41));
    defparam i3_4_lut_adj_67.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_68 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n601));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_68.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_69 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n592));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_69.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_70 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n598));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_70.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_71 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n589));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_71.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_72 (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n628));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_72.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_73 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[10]), .O(n32));
    defparam i3_4_lut_adj_73.LUT_INIT = 16'h0400;
    SB_LUT4 i13171_2_lut_3_lut (.I0(\preSatVoltage[21] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[12] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13171_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i13169_2_lut_3_lut (.I0(\preSatVoltage[19] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[10] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13169_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_74 (.I0(\preSatVoltage[19] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n538));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_74.LUT_INIT = 16'h00d0;
    SB_LUT4 i3_4_lut_adj_75 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[9]), .O(n29));
    defparam i3_4_lut_adj_75.LUT_INIT = 16'h0400;
    SB_LUT4 i3_4_lut_adj_76 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[5]), .O(n17));
    defparam i3_4_lut_adj_76.LUT_INIT = 16'h0400;
    SB_LUT4 D_15__I_0_10_i49_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[7]), .O(n71));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i49_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i57_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[11]), .O(n83));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i57_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i41_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[3]), .O(n59));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i41_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i35_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[0]), .O(n50));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i35_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i63_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[14]), .O(n92));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i63_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i47_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[6]), .O(n68));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i47_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i43_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[4]), .O(n62));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i43_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i37_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[1]), .O(n53));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i37_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i45_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[5]), .O(n65));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i45_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_adj_77 (.I0(Out_31__N_332), .I1(\preSatVoltage[9] ), 
            .I2(Out_31__N_333), .I3(Look_Up_Table_out1_1[12]), .O(n38));
    defparam i3_4_lut_adj_77.LUT_INIT = 16'h0400;
    SB_LUT4 D_15__I_0_10_i39_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[2]), .O(n56));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i39_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i55_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[10]), .O(n80));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i55_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_78 (.I0(\preSatVoltage[13] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n244));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_78.LUT_INIT = 16'h00d0;
    SB_LUT4 D_15__I_0_10_i158_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), 
            .O(n233));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i158_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 equal_13243_i14_2_lut_3_lut_3_lut (.I0(\preSatVoltage[13] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(n14_adj_6));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam equal_13243_i14_2_lut_3_lut_3_lut.LUT_INIT = 16'h5858;
    SB_LUT4 D_15__I_0_10_i136_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), 
            .O(n200));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i136_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i138_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), 
            .O(n203));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i138_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_i39_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(\Product_mul_temp[26] ), .O(n86));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_i39_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i53_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[9]), .O(n77));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i53_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i134_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), 
            .O(n197));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i134_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i162_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), 
            .O(n239));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i162_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i140_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), 
            .O(n206));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i140_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i59_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[12]), .O(n86_adj_7));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i59_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i146_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[6]), .I3(Out_31__N_332), 
            .O(n215));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i146_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i61_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[13]), .O(n89));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i61_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i51_2_lut_4_lut (.I0(Out_31__N_332), .I1(Out_31__N_333), 
            .I2(\preSatVoltage[10] ), .I3(Look_Up_Table_out1_1[8]), .O(n74));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam D_15__I_0_10_i51_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 D_15__I_0_10_i154_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), 
            .O(n227));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i154_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_i138_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), .I1(Out_31__N_333), 
            .I2(\Product_mul_temp[26] ), .I3(Out_31__N_332), .O(n233_adj_8));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_i138_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i152_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), 
            .O(n224));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i152_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i150_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[8]), .I3(Out_31__N_332), 
            .O(n221));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i150_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i142_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), 
            .O(n209));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i142_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i160_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), 
            .O(n236));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i160_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i156_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), 
            .O(n230));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i156_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_79 (.I0(\preSatVoltage[13] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n244_adj_9));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_79.LUT_INIT = 16'h00d0;
    SB_LUT4 D_15__I_0_10_i144_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), 
            .O(n212));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i144_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 D_15__I_0_10_i148_2_lut_3_lut_4_lut (.I0(\preSatVoltage[13] ), 
            .I1(Out_31__N_333), .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), 
            .O(n218));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam D_15__I_0_10_i148_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_80 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n279));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_80.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_81 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[8]), .I3(Out_31__N_332), .O(n270));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_81.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_82 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), .O(n267));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_82.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_83 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n255));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_83.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_84 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n285));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_84.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_85 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[6]), .I3(Out_31__N_332), .O(n264));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_85.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_86 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n258));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_86.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_87 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n249));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_87.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_88 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n246));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_88.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_89 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), .O(n273));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_89.LUT_INIT = 16'h00e0;
    SB_LUT4 i13173_2_lut_3_lut (.I0(\preSatVoltage[23] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[14] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13173_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_90 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), .O(n282));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_90.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_91 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n261));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_91.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_92 (.I0(\preSatVoltage[23] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n19681));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_92.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_93 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), .O(n288));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_93.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_94 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), .O(n276));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_94.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_95 (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n252));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_95.LUT_INIT = 16'h00e0;
    SB_LUT4 i13164_2_lut_3_lut (.I0(\preSatVoltage[14] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[5] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13164_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_3_lut_4_lut (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[13]), .I3(Out_31__N_332), .O(n789));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_96 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[12]), .I3(Out_31__N_332), .O(n785));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_96.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_97 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[7]), .I3(Out_31__N_332), .O(n765));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_97.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_98 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[4]), .I3(Out_31__N_332), .O(n753));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_98.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_99 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[1]), .I3(Out_31__N_332), .O(n741));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_99.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_100 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[5]), .I3(Out_31__N_332), .O(n757));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_100.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_101 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[2]), .I3(Out_31__N_332), .O(n745));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_101.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_102 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[6]), .I3(Out_31__N_332), .O(n761));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_102.LUT_INIT = 16'h000e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_103 (.I0(\preSatVoltage[12] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[15]), .I3(Out_31__N_332), .O(n195));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_2_lut_3_lut_4_lut_adj_103.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_3_lut_4_lut_adj_104 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[0]), .I3(Out_31__N_332), .O(n737));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_104.LUT_INIT = 16'h000e;
    SB_LUT4 i13162_2_lut_3_lut (.I0(\preSatVoltage[12] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[3] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13162_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_3_lut_4_lut_adj_105 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[3]), .I3(Out_31__N_332), .O(n749));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_105.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_106 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[11]), .I3(Out_31__N_332), .O(n781));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_106.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_107 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[10]), .I3(Out_31__N_332), .O(n777));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_107.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_108 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[9]), .I3(Out_31__N_332), .O(n773));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_108.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_109 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[8]), .I3(Out_31__N_332), .O(n769));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_109.LUT_INIT = 16'h000e;
    SB_LUT4 i1_3_lut_4_lut_adj_110 (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Look_Up_Table_out1_1[14]), .I3(Out_31__N_332), .O(n19684));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i1_3_lut_4_lut_adj_110.LUT_INIT = 16'h000e;
    SB_LUT4 i13174_2_lut_3_lut (.I0(\preSatVoltage[24] ), .I1(Out_31__N_333), 
            .I2(Out_31__N_332), .I3(GND_net), .O(\dVoltage[15] ));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(52[15] 53[18])
    defparam i13174_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_111 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[14]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n435));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_111.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_112 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[14]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n141));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_112.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_113 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[14]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n631));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_113.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_114 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[6]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[11] ), .O(n117));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_114.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_115 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[6]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[17] ), .O(n411));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_115.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_116 (.I0(Out_31__N_332), .I1(Look_Up_Table_out1_1[6]), 
            .I2(Out_31__N_333), .I3(\preSatVoltage[21] ), .O(n607));   // ../../hdlcoderFocCurrentFixptHdl/Saturate_Output.v(51[36] 53[19])
    defparam i1_2_lut_3_lut_4_lut_adj_116.LUT_INIT = 16'h4440;
    
endmodule
