// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sat Jun  1 16:19:04 2019
//
// Verilog Description of module DarkRoomOOTXdecoder
//

module DarkRoomOOTXdecoder (clock, reset, address, read, readdata, 
            write, writedata, waitrequest, uart_tx, sensor_signals, 
            led) /* synthesis syn_module_defined=1 */ ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(39[8:27])
    input clock;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(40[8:13])
    input reset;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(41[8:13])
    input [5:0]address;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    input read;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(44[8:12])
    output [31:0]readdata;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(45[23:31])
    input write;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(46[8:13])
    input [31:0]writedata;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(47[22:31])
    output waitrequest;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(48[9:20])
    output uart_tx;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(50[9:16])
    input [7:0]sensor_signals;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(51[32:46])
    output [7:0]led;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(52[15:18])
    
    wire clock_c /* synthesis SET_AS_NETWORK=clock_c, is_clock=1 */ ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(40[8:13])
    
    wire GND_net, VCC_net, reset_c, address_c_5, address_c_4, address_c_3, 
        address_c_2, address_c_1, address_c_0, readdata_c_31, readdata_c_30, 
        readdata_c_29, readdata_c_28, readdata_c_27, readdata_c_26, 
        readdata_c_25, readdata_c_24, readdata_c_23, readdata_c_22, 
        readdata_c_21, readdata_c_20, readdata_c_19, readdata_c_18, 
        readdata_c_17, readdata_c_16, readdata_c_15, readdata_c_14, 
        readdata_c_13, readdata_c_12, readdata_c_11, readdata_c_10, 
        readdata_c_9, readdata_c_8, readdata_c_7, readdata_c_6, readdata_c_5, 
        readdata_c_4, readdata_c_3, readdata_c_2, readdata_c_1, readdata_c_0, 
        write_c, writedata_c_31, writedata_c_30, writedata_c_29, writedata_c_28, 
        writedata_c_27, writedata_c_26, writedata_c_25, writedata_c_24, 
        writedata_c_23, writedata_c_22, writedata_c_21, writedata_c_20, 
        writedata_c_19, writedata_c_18, writedata_c_17, writedata_c_16, 
        writedata_c_15, writedata_c_14, writedata_c_13, writedata_c_12, 
        writedata_c_11, writedata_c_10, writedata_c_9, writedata_c_8, 
        writedata_c_7, writedata_c_6, writedata_c_5, writedata_c_4, 
        writedata_c_3, writedata_c_2, writedata_c_1, writedata_c_0, 
        waitrequest_c, sensor_signals_c_7, sensor_signals_c_6, sensor_signals_c_5, 
        sensor_signals_c_4, sensor_signals_c_3, sensor_signals_c_2, sensor_signals_c_1, 
        sensor_signals_c_0, led_c_7, led_c_6, led_c_5, led_c_4, led_c_3, 
        led_c_2, led_c_1, led_c_0;
    wire [31:0]sensor_select;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(98[12:25])
    wire [1:0]sync;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(116[12:16])
    wire [271:0]n4568;
    wire [271:0]n4551;
    wire [31:0]\ootx_crc32_o[1] ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(119[13:25])
    wire [31:0]\ootx_crc32_o[0] ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(119[13:25])
    
    wire n524, n525, n37, n8, n1032, n1030, n1028, n1026, n1024, 
        n1022, n1020, n1018, n1016, n1014, n1012, n1010, n1008, 
        n1006, n1004, n1002, n1000, n998, n996, n994, n992, 
        n990, n988, n986, n984, n982, n980, n978, n976, n974, 
        n972, n970, n968, n966, n964, n962, n960, n958, n956, 
        n954, n952, n950, n948, n946, n944, n942, n940, n938, 
        n936, n934, n932, n930, n928, n926, n924, n922, n920, 
        n918, n916, n914, n912, n910, n908, n906, n904, n902, 
        n900, n898, n896, n894, n892, n890, n888, n886, n884, 
        n882, n880, n878, n876, n874, n872, n870, n868, n866, 
        n864, n862, n860, n858, n856, n854, n852, n850, n848, 
        n846, n844, n842, n840, n838, n836, n834, n832, n830, 
        n828, n826, n824, n822, n820, n818, n816, n814, n812, 
        n810, n808, n806, n804, n802, n800, n798, n796, n794, 
        n792, n790, n788, n786, n784, n782, n780, n778, n776, 
        n774, n772, n770, n768, n766, n764, n762, n760, n758, 
        n756, n754, n752, n750, n748, n746, n744, n742, n740, 
        n738, n736, n734, n732, n730, n728, n726, n724, n722, 
        n720, n718, n716, n714, n712, n710, n708, n706, sensor_N_132, 
        sensor_state;
    wire [31:0]counter_from_last_rise;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    
    wire data;
    wire [1:0]\ootx_states[1] ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(52[9:20])
    wire [1:0]\ootx_states[0] ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(52[9:20])
    
    wire new_data;
    wire [30:0]lighthouse;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(60[9:19])
    
    wire n704, n702, n4099, n4100, n4101, n4102, n4103, n4104, 
        n4105, n24315;
    wire [1:0]ootx_payloads_N_1744;
    
    wire n45, n338, n339, n340, n341, n342, n343, n344, n345, 
        n346, n347, n348, n349, n350, n351, n352, n353, n354, 
        n355, n356, n357, n358, n359, n360, n361, n362, n363, 
        n364, n365, n366, n367, n368;
    wire [15:0]ootx_payloads_N_1730;
    
    wire ootx_payloads_N_1698, n1170, n1171, n1172, n1173, n1174, 
        n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
        n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
        n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
        n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
        n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
        n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
        n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
        n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
        n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
        n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
        n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
        n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
        n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
        n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
        n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
        n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
        n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
        n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
        n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
        n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
        n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
        n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
        n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
        n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
        n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
        n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
        n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
        n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
        n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
        n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
        n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
        n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
        n1431, n1432, n1433, n23005, n23007, n23009, n23011, n23013, 
        n23015, n23017, n23019, n23021, n23023, n23025, n23027, 
        n23029, n23031, n23033, n23035, n23037, n23039, n23041, 
        n23043, n23045, n23047, n23049, n23051, n23053, n23055, 
        n23057, n23059, n23061, n23063, n23065, n23067, n23069, 
        n23071, n23001, n23073, n23075, n23077, n23079, n23081, 
        n23083, n23085, n23087, n23089, n23091, n23093, n23095, 
        n23097, n23099, n23101, n23103, n23105, n23107, n23109, 
        n23111, n23113, n23115, n23117, n23119, n23121, n23123, 
        n23125, n23477, n23479, n23481, n23483, n23485, n23487, 
        n23489, n23491, n23493, n23495, n23497, n23499, n23501, 
        n23503, n23505, n23507, n23509, n23511, n23471, n23465, 
        n23459, n23453, n23447, n23441, n23435, n23429, n23423, 
        n23417, n23411, n23401, n23391, n23513, n23515, n23517, 
        n23519, n23521, n23523, n23525, n23527, n23529, n23531, 
        n23533, n23535, n23537, n23539, n23541, n23543, n23545, 
        n1, n23641, n25888, n4673, n30, n28, n26, n24, n22, 
        n20, n18, n16, n2852, n2853, n2854, n2855, n2856, n2857, 
        n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, 
        n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
        n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
        n2882;
    wire [30:0]ootx_payloads_N_1699;
    
    wire n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
        n3088, n3089, n3090, n3091, n3092, n3093_adj_2243, n3094_adj_2244, 
        n3095_adj_2245, n3096_adj_2246, n3097_adj_2247, n3098_adj_2248, 
        n3099_adj_2249, n3100_adj_2250, n3101, n3102, n3103, n3104, 
        n3105, n3106, n3107, n3108, n3109, n3110, n3111, n14, 
        n12, n10, n4702, n4700, n23475, n23469, n8_adj_2251, n588, 
        n590, n592, n594, n596, n20_adj_2252, n700, n698, n696, 
        n694, n692, n690, n23463, n23457, n23451, n23445, n23439, 
        n23433, n23427, n23421, n23415, n23409, n23399, n12201, 
        n12200, n12199, n12198, n12197, n12196, n12195, n12194, 
        n12193, n12192, n12191, n12190, n12189, n12188, n12187, 
        n12186, n12185, n12184, n12183, n12182, n12181, n12180, 
        n12179, n12178, n12177, n12176, n12175, n12174, n12173, 
        n12172, n12171, n12170, n12169, n12168, n12167, n12166, 
        n12165, n12164, n12163, n12162, n12161, n12160, n12159, 
        n12158, n12157, n12156, n12155, n12154, n12153, n12152, 
        n12151, n12150, n12149, n12148, n12147, n12146, n12145, 
        n12144, n12143, n12142, n12141, n12140, n12139, n12138, 
        n12137, n12136, n12135, n12134, n12133, n12132, n12131, 
        n12130, n12129, n12128, n12127, n12126, n12125, n12124, 
        n12123, n12122, n12121, n12120, n12119, n12118, n12117, 
        n12116, n12115, n12114, n12113, n12112, n12111, n12110, 
        n12109, n12108, n12107, n12106, n12105, n12104, n12103, 
        n12102, n12101, n12100, n12099, n12098, n12097, n12096, 
        n12095, n12094, n12093, n12092, n12091, n12090, n12089, 
        n12088, n12087, n12086, n12085, n12084, n12083, n12082, 
        n12081, n12080, n12079, n12078, n12077, n12076, n12075, 
        n12074, n12073, n12072, n12071, n12070, n12069, n12068, 
        n12067, n12066, n12065, n12064, n12063, n12062, n12061, 
        n12060, n12059, n12058, n12057, n12056, n12055, n12054, 
        n12053, n12052, n12051, n12050, n12049, n12048, n12047, 
        n12046, n12045, n12044, n12043, n12042, n12041, n12040, 
        n12039, n12038, n12037, n12036, n12035, n12034, n12033, 
        n12032, n12031, n12030, n12029, n12028, n12027, n12026, 
        n12025, n12024, n12023, n12022, n12021, n12020, n12019, 
        n12018, n12017, n12016, n12015, n12014, n12013, n12012, 
        n12011, n12010, n12009, n12008, n12007, n12006, n12005, 
        n12004, n12003, n12002, n12001, n12000, n11999, n11998, 
        n11997, n11996, n11995, n11994, n11993, n11992, n11991, 
        n11990, n11989, n11988, n11987, n11986, n11985, n11984, 
        n11983, n11982, n11981, n11980, n11979, n11978, n11977, 
        n11976, n11975, n11974, n11973, n11972, n11971, n11970, 
        n11969, n11968, n11967, n11966, n11965, n11964, n11963, 
        n11962, n11961, n11960, n11959, n11958, n11957, n11956, 
        n11955, n11954, n11953, n36, n35, n17, n24248, n24245, 
        n24242, n24239, n24236, n24233, payload_lengths_1_0, payload_lengths_0_0, 
        n11952, n11951, n11950, n11949, n11948, n11947, n11946, 
        n11945, n11944, n11943, n11942, n11941, n11940, n11939, 
        n13329, crc32s_1_31, crc32s_1_30, crc32s_1_29, crc32s_1_28, 
        crc32s_1_27, crc32s_1_26, crc32s_1_25, crc32s_1_24, crc32s_1_23, 
        crc32s_1_22, crc32s_1_21, crc32s_1_20, crc32s_1_19, crc32s_1_18, 
        crc32s_1_17, crc32s_1_16, crc32s_1_15, crc32s_1_14, crc32s_1_13, 
        crc32s_1_12, crc32s_1_11, crc32s_1_10, crc32s_1_9, crc32s_1_8, 
        crc32s_1_7, crc32s_1_6, crc32s_1_5, crc32s_1_4, crc32s_1_3, 
        crc32s_1_2, crc32s_1_1, crc32s_1_0, n11612, n11611, n11610, 
        n11609, n11608, n11607, n11606, n11605, n11604, n11602, 
        n23003, n11600, n11599, n11598, n11597, n11596, n11595, 
        n11594, n11593, n11592, n11591, n11590, n11589, n11588, 
        n11587, n11586, n11585, n11584, n11583, n11582, n11581, 
        n11580, n11579, n11578, n11577, n11576, n11575, n11574, 
        n11573, n11572, n11571, n11570, n11569, n11568, n11567, 
        n11566, n11565, n11564, n11563, n11562, n11561, n11560, 
        n11559, n11558, n11557, n11556, n11555, n11554, n11553, 
        n11552, n11551, n11550, n11549, n11548, n11547, n11546, 
        n11545, n11544, n11543, n11542, n11541, n11540, n11539, 
        n11538, n11537, n11536, n11535, n11534, n11533, n11532, 
        n11531, n11530, n11529, n11528, n11527, n11526, n11525, 
        n11524, n11523, n11522, n11521, n11520, n11519, n11518, 
        n11517, n11516, n11515, n11514, n11513, n11512, n11511, 
        n11510, n11509, n11508, n11507, n11506, n11505, n11504, 
        n11503, n11502, n11501, n11500, n11499, n11498, n11497, 
        n11496, n11495, n11494, n11493, n11492, n11491, n11490, 
        n11489, n11488, n11487, n11486, n11485, n11484, n11483, 
        n11482, n11481, n11480, n11479, n11478, n11477, n11476, 
        n11475, n11474, n11473, n11472, n11471, n11470, n11469, 
        n11468, n11467, n11466, n11465, n11464, n11463, n11462, 
        n11461, n11460, n11459, n11458, n11457, n11456, n11455, 
        n11454, n11453, n11452, n11451, n11450, n11449, n11448, 
        n11447, n11446, n11445, n11444, n11443, n11442, n11441, 
        n11440, n11439, n11438, n11437, n11436, n11435, n11434, 
        n11433, n11432, n11431, n11430, n11429, n11428, n11427, 
        n11426, n11425, n11424, n11423, n11422, n11421, n11420, 
        n11419, n11418, n11417, n11416, n11415, n11414, n11413, 
        n11412, n11411, n11410, n11409, n11408, n11407, n11406, 
        n11405, n11404, n11403, n11402, n11401, n11400, n11399, 
        n11398, n11397, n11396, n11395, n11394, n11393, n11392, 
        n11391, n11390, n11389, n11388, n11387, n11386, n11385, 
        n11384, n11383, n11382, n11381, n11380, n11379, n11378, 
        n11377, n11376, n11375, n11374, n11373, n11372, n11371, 
        n11370, n11369, n11368, n11367, n11366, n11365, n523, 
        n11364, n11363, n11362, n11361, n11360, n11359, n11358, 
        n11357, n11356, n72, n24282, n24306, n3917, n3916, n3915, 
        n3913, n3912, n11355, n8_adj_2253, n8_adj_2254, n8_adj_2255, 
        n1_adj_2256, n24522, n24468, n11354, n11353, n11352, n11351, 
        n11350, n24152, n11349, n688, n686, n684, n682, n680, 
        n11348, n678, n676, n674, n672, n670, n668, n666, n664, 
        n662, n660, n658, n656, n654, n652, n650, n648, n646, 
        n644, n642, n640, n638, n636, n634, n632, n630, n628, 
        n626, n624, n622, n620, n618, n616, n614, n11347, n11346, 
        n11345, n11344, n11343, n11342, n11341, n11340, n35_adj_2257, 
        n11339, n11338, n11337, n11336, n11335, n11334, n11333, 
        n13221, n11332, n2680, n11331, n11330, n11329, n11328, 
        n2282, n11327, n527, n11326, n11325, n9797, n11324, n11323, 
        n3805, n11322, n3804, n11321, n3803, n3802, n3801, n3800, 
        n11320, n3799, n11319, n11318, n2208, n24501, n11317, 
        n11316, n11315, n11314, n11313, n598, n600, n602, n608, 
        n606, n11312, n11311, n11310, n9771, n11309, n3737, n3736, 
        n3735, n3734, n3733, n3732, n3731, n3730, n3729, n3728, 
        n3727, n3726, n3725, n3724, n3723, n24453, n3696, n3695, 
        n3694, n3693, n3692, n3691, n3690, n3689, n11308, n24417, 
        n11307, n586, n11306, n11305, n580, n11304, n584, n24525, 
        n24465, n24528, n24462, n24531, n24459, n582, n11303, 
        n11302, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
        n4303, n24393, n576, n574, n572, n570, n568, n566, n11301, 
        n11300, n24534, n24456, n24363, n24519, n4, n526, n11299, 
        n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, 
        n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
        n11298, n11297, n11296, n11295, n11294, n11293, n11292, 
        n11291, n529, n24516, n11290, n24513, n542, n540, n556, 
        n11289, n11288, n554, n4218, n4219, n4220, n4221, n4222, 
        n4223, n4224, n4225, n11287, n521, n11286, n11285, n6334, 
        n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, 
        n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, 
        n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, 
        n6359, n6361, n6362, n6363, n6364, n6365, n564, n562, 
        n560, n612, n4237, n4238, n4239, n4240, n4241, n4242, 
        n4243, n4244, n24498, n24366, n24495, n3100, n3099, n3098, 
        n3097, n3096, n3095, n3094, n3093, n2679, n610, n558, 
        n578, n19468, n8_adj_2258, n24147, n54, n8_adj_2259, n530, 
        n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, 
        n552, n550, n548, data_N_1808, n546, n544, n24309, n8_adj_2260, 
        n24492, n4090, n528, n4091, n4092, n604, n533, n532, 
        n531, n4150, n4093, n4094, n4095, n4151, n4152, n4153, 
        n4154, n4155, n4156, n4157, n4096, n538, n536, n535, 
        n534, n8_adj_2261, n24507, n2, n24489, n8_adj_2262, n23974, 
        n4097, n24312, n8_adj_2263, n24504, n4098, ootx_payloads_1_263, 
        ootx_payloads_1_262, ootx_payloads_1_261, ootx_payloads_1_260, 
        ootx_payloads_1_259, ootx_payloads_1_258, ootx_payloads_1_257, 
        ootx_payloads_1_256, ootx_payloads_1_255, ootx_payloads_1_254, 
        ootx_payloads_1_253, ootx_payloads_1_252, ootx_payloads_1_251, 
        ootx_payloads_1_250, ootx_payloads_1_249, ootx_payloads_1_248, 
        ootx_payloads_1_247, ootx_payloads_1_246, ootx_payloads_1_245, 
        ootx_payloads_1_244, ootx_payloads_1_243, ootx_payloads_1_242, 
        ootx_payloads_1_241, ootx_payloads_1_240, ootx_payloads_1_239, 
        ootx_payloads_1_238, ootx_payloads_1_237, ootx_payloads_1_236, 
        ootx_payloads_1_235, ootx_payloads_1_234, ootx_payloads_1_233, 
        ootx_payloads_1_232, ootx_payloads_1_231, ootx_payloads_1_230, 
        ootx_payloads_1_229, ootx_payloads_1_228, ootx_payloads_1_227, 
        ootx_payloads_1_226, ootx_payloads_1_225, ootx_payloads_1_224, 
        ootx_payloads_1_223, ootx_payloads_1_222, ootx_payloads_1_221, 
        ootx_payloads_1_220, ootx_payloads_1_219, ootx_payloads_1_218, 
        ootx_payloads_1_217, ootx_payloads_1_216, ootx_payloads_1_215, 
        ootx_payloads_1_214, ootx_payloads_1_213, ootx_payloads_1_212, 
        ootx_payloads_1_211, ootx_payloads_1_210, ootx_payloads_1_209, 
        ootx_payloads_1_208, ootx_payloads_1_207, ootx_payloads_1_206, 
        ootx_payloads_1_205, ootx_payloads_1_204, ootx_payloads_1_203, 
        ootx_payloads_1_202, ootx_payloads_1_201, ootx_payloads_1_200, 
        ootx_payloads_1_199, ootx_payloads_1_198, ootx_payloads_1_197, 
        ootx_payloads_1_196, ootx_payloads_1_195, ootx_payloads_1_194, 
        ootx_payloads_1_193, ootx_payloads_1_192, ootx_payloads_1_191, 
        ootx_payloads_1_190, ootx_payloads_1_189, ootx_payloads_1_188, 
        ootx_payloads_1_187, ootx_payloads_1_186, ootx_payloads_1_185, 
        ootx_payloads_1_184, ootx_payloads_1_183, ootx_payloads_1_182, 
        ootx_payloads_1_181, ootx_payloads_1_180, ootx_payloads_1_179, 
        ootx_payloads_1_178, ootx_payloads_1_177, ootx_payloads_1_176, 
        ootx_payloads_1_175, ootx_payloads_1_174, ootx_payloads_1_173, 
        ootx_payloads_1_172, ootx_payloads_1_171, ootx_payloads_1_170, 
        ootx_payloads_1_169, ootx_payloads_1_168, ootx_payloads_1_167, 
        ootx_payloads_1_166, ootx_payloads_1_165, ootx_payloads_1_164, 
        ootx_payloads_1_163, ootx_payloads_1_162, ootx_payloads_1_161, 
        ootx_payloads_1_160, ootx_payloads_1_159, ootx_payloads_1_158, 
        ootx_payloads_1_157, ootx_payloads_1_156, ootx_payloads_1_155, 
        ootx_payloads_1_154, ootx_payloads_1_153, ootx_payloads_1_152, 
        ootx_payloads_1_151, ootx_payloads_1_150, ootx_payloads_1_149, 
        ootx_payloads_1_148, ootx_payloads_1_147, ootx_payloads_1_146, 
        ootx_payloads_1_145, ootx_payloads_1_144, ootx_payloads_1_143, 
        ootx_payloads_1_142, ootx_payloads_1_141, ootx_payloads_1_140, 
        ootx_payloads_1_139, ootx_payloads_1_138, ootx_payloads_1_137, 
        ootx_payloads_1_136, ootx_payloads_1_135, ootx_payloads_1_134, 
        ootx_payloads_1_133, ootx_payloads_1_132, ootx_payloads_1_131, 
        ootx_payloads_1_130, ootx_payloads_1_129, ootx_payloads_1_128, 
        ootx_payloads_1_127, ootx_payloads_1_126, ootx_payloads_1_125, 
        ootx_payloads_1_124, ootx_payloads_1_123, ootx_payloads_1_122, 
        ootx_payloads_1_121, ootx_payloads_1_120, ootx_payloads_1_119, 
        ootx_payloads_1_118, ootx_payloads_1_117, ootx_payloads_1_116, 
        ootx_payloads_1_115, ootx_payloads_1_114, ootx_payloads_1_113, 
        ootx_payloads_1_112, ootx_payloads_1_111, ootx_payloads_1_110, 
        ootx_payloads_1_109, ootx_payloads_1_108, ootx_payloads_1_107, 
        ootx_payloads_1_106, ootx_payloads_1_105, ootx_payloads_1_104, 
        ootx_payloads_1_103, ootx_payloads_1_102, ootx_payloads_1_101, 
        ootx_payloads_1_100, ootx_payloads_1_99, ootx_payloads_1_98, ootx_payloads_1_97, 
        ootx_payloads_1_96, ootx_payloads_1_95, ootx_payloads_1_94, ootx_payloads_1_93, 
        ootx_payloads_1_92, ootx_payloads_1_91, ootx_payloads_1_90, ootx_payloads_1_89, 
        ootx_payloads_1_88, ootx_payloads_1_87, ootx_payloads_1_86, ootx_payloads_1_85, 
        ootx_payloads_1_84, ootx_payloads_1_83, ootx_payloads_1_82, ootx_payloads_1_81, 
        ootx_payloads_1_80, ootx_payloads_1_79, ootx_payloads_1_78, ootx_payloads_1_77, 
        ootx_payloads_1_76, ootx_payloads_1_75, ootx_payloads_1_74, ootx_payloads_1_73, 
        ootx_payloads_1_72, ootx_payloads_1_71, ootx_payloads_1_70, ootx_payloads_1_69, 
        ootx_payloads_1_68, ootx_payloads_1_67, ootx_payloads_1_66, ootx_payloads_1_65, 
        ootx_payloads_1_64, ootx_payloads_1_63, ootx_payloads_1_62, ootx_payloads_1_61, 
        ootx_payloads_1_60, ootx_payloads_1_59, ootx_payloads_1_58, ootx_payloads_1_57, 
        ootx_payloads_1_56, ootx_payloads_1_55, ootx_payloads_1_54, ootx_payloads_1_53, 
        ootx_payloads_1_52, ootx_payloads_1_51, ootx_payloads_1_50, ootx_payloads_1_49, 
        ootx_payloads_1_48, ootx_payloads_1_47, ootx_payloads_1_46, ootx_payloads_1_45, 
        ootx_payloads_1_44, ootx_payloads_1_43, ootx_payloads_1_42, ootx_payloads_1_41, 
        ootx_payloads_1_40, ootx_payloads_1_39, ootx_payloads_1_38, ootx_payloads_1_37, 
        ootx_payloads_1_36, ootx_payloads_1_35, ootx_payloads_1_34, ootx_payloads_1_33, 
        ootx_payloads_1_32, ootx_payloads_1_31, ootx_payloads_1_30, ootx_payloads_1_29, 
        ootx_payloads_1_28, ootx_payloads_1_27, ootx_payloads_1_26, ootx_payloads_1_25, 
        ootx_payloads_1_24, ootx_payloads_1_23, ootx_payloads_1_22, ootx_payloads_1_21, 
        ootx_payloads_1_20, ootx_payloads_1_19, ootx_payloads_1_18, ootx_payloads_1_17, 
        ootx_payloads_1_16, ootx_payloads_1_15, ootx_payloads_1_14, ootx_payloads_1_13, 
        ootx_payloads_1_12, ootx_payloads_1_11, ootx_payloads_1_10, ootx_payloads_1_9, 
        ootx_payloads_1_8, ootx_payloads_1_7, ootx_payloads_1_6, ootx_payloads_1_5, 
        ootx_payloads_1_4, ootx_payloads_1_3, ootx_payloads_1_2, ootx_payloads_1_1, 
        ootx_payloads_1_0, n522, n8917, n24833, n24832, n24831, 
        n24830, n24826, n24825, n8_adj_2264, n24030, n8_adj_2265, 
        n24815, n24814, n8_adj_2266, n24812, n23639, n24801, n24800, 
        n24799, n24798, n24797, n24796, n24795, n24794, n4671, 
        n24783, data_counters_0_0, data_counters_0_1, data_counters_0_2, 
        data_counters_0_3, data_counters_0_4, data_counters_0_5, data_counters_0_6, 
        data_counters_0_7, data_counters_0_8, data_counters_0_9, data_counters_0_10, 
        data_counters_0_11, data_counters_0_12, data_counters_0_13, data_counters_0_14, 
        data_counters_0_15, data_counters_0_16, data_counters_0_17, data_counters_0_18, 
        data_counters_0_19, data_counters_0_20, data_counters_0_21, data_counters_0_22, 
        data_counters_0_23, data_counters_0_24, data_counters_0_25, data_counters_0_26, 
        data_counters_0_27, data_counters_0_28, data_counters_0_29, data_counters_0_30, 
        data_counters_1_0, data_counters_1_1, data_counters_1_2, data_counters_1_3, 
        data_counters_1_4, data_counters_1_5, data_counters_1_6, data_counters_1_7, 
        data_counters_1_8, data_counters_1_9, data_counters_1_10, data_counters_1_11, 
        data_counters_1_12, data_counters_1_13, data_counters_1_14, data_counters_1_15, 
        data_counters_1_16, data_counters_1_17, data_counters_1_18, data_counters_1_19, 
        data_counters_1_20, data_counters_1_21, data_counters_1_22, data_counters_1_23, 
        data_counters_1_24, data_counters_1_25, data_counters_1_26, data_counters_1_27, 
        data_counters_1_28, data_counters_1_29, data_counters_1_30, bit_counters_0_0, 
        bit_counters_0_1, bit_counters_0_2, bit_counters_0_3, bit_counters_0_4, 
        bit_counters_0_5, bit_counters_0_6, bit_counters_0_7, bit_counters_0_8, 
        bit_counters_0_9, bit_counters_0_10, bit_counters_0_11, bit_counters_0_12, 
        bit_counters_0_13, bit_counters_0_14, bit_counters_0_15, bit_counters_0_16, 
        bit_counters_0_17, bit_counters_0_18, bit_counters_0_19, bit_counters_0_20, 
        bit_counters_0_21, bit_counters_0_22, bit_counters_0_23, bit_counters_0_24, 
        bit_counters_0_25, bit_counters_0_26, bit_counters_0_27, bit_counters_0_28, 
        bit_counters_0_29, bit_counters_0_30, bit_counters_1_0, bit_counters_1_1, 
        bit_counters_1_2, bit_counters_1_3, bit_counters_1_4, bit_counters_1_5, 
        bit_counters_1_6, bit_counters_1_7, bit_counters_1_8, bit_counters_1_9, 
        bit_counters_1_10, bit_counters_1_11, bit_counters_1_12, bit_counters_1_13, 
        bit_counters_1_14, bit_counters_1_15, bit_counters_1_16, bit_counters_1_17, 
        bit_counters_1_18, bit_counters_1_19, bit_counters_1_20, bit_counters_1_21, 
        bit_counters_1_22, bit_counters_1_23, bit_counters_1_24, bit_counters_1_25, 
        bit_counters_1_26, bit_counters_1_27, bit_counters_1_28, bit_counters_1_29, 
        bit_counters_1_30, n11016, n24782, n24781, n25885, n25882, 
        n25879, n25876, n25873, n25870, n25867, n25864, n25861, 
        n1_adj_2267, n25858, n25855, n25852, n25849, n25846, n25843, 
        n25840, n25837, n25831, n8_adj_2268, n25825, n25822, n25819, 
        n25816, n25813, n25810, n25807, n25804, n25801, n25798, 
        n25795, n25792, n25789, n25783, n25777, n25774, n25771, 
        n25768, n25765, n25762, n24018, n25759, n25756, n25753, 
        n25750, n25747, n25744, n25741, n25738, n25735, n25732, 
        n25729, n25726, n25723, n25717, n25711, n25705, n25699, 
        n25693, n25687, n25681, n25675, n25669, n25663, n25657, 
        n25651, n25645, n25639, n25636, n25633, n25630, n25627, 
        n25624, n25621, n25615, n25612, n25609, n25606, n25603, 
        n25597, n24780, n25594, n25591, n25588, n25585, n25579, 
        n25576, n25573, n25570, n25567, n25564, n8_adj_2269, n24779, 
        n25561, n25558, n25555, n25552, n25549, n25543, n25540, 
        n25537, n25531, n24778, n24777, n24776, n25525, n25519, 
        n25513, n25507, n25501, n25495, n24775, n24774, n25489, 
        n25483, n25477, n25471, n25465, n25462, n25459, n25456, 
        n24773, n24486, n25453, n25447, n25441, n25435, n25429, 
        n25423, n25417, n24772, n24771, n24770, n24769, n24768, 
        n24767, n24765, n25411, n25405, n25402, n25399, n25396, 
        n25393, n25390, n25387, n25381, n25378, n24763, n24761, 
        n24759, n25375, n25372, n25369, n25366, n25363, n25360, 
        n25357, n25354, n25351, n25348, n25345, n25339, n25336, 
        n25333, n25330, n25327, n25324, n25321, n25318, n25315, 
        n25312, n25309, n25306, n25303, n25297, n25291, n25285, 
        n25279, n25273, n25267, n25264, n25261, n25258, n25255, 
        n25252, n25249, n25246, n25243, n25240, n25237, n25234, 
        n25231, n25228, n25225, n25216, n25213, n25210, n25207, 
        n25204, n25201, n9200, n23971, n22997, n24731, n37_adj_2270, 
        n38, n39, n40, n41, n42, n43, n44, n45_adj_2271, n46, 
        n47, n48, n49, n50, n51, n52, n53, n54_adj_2272, n55, 
        n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
        n66, n67, n68, n24730, n24729, n24728, n24727, n24726, 
        n24725, n24724, n8_adj_2273, n8_adj_2274, n23407, n24692, 
        n8_adj_2275, n28_adj_2276, n8_adj_2277, n23397, n8_adj_2278, 
        n23972, n24666, n8_adj_2279, n24665, n24664, n24663, n24662, 
        n24661, n24660, n24659, n24658, n24657, n24656, n24655, 
        n24654, n24653, n8_adj_2280, n23389, n24643, n24642, n24639, 
        n24635, n24634, n24628, n24627, n24626, n24625, n24624, 
        n24623, n24622, n24620, n24617, n24616, n29, n8_adj_2281, 
        n23697, n8_adj_2282, n33, n13397, n13402, n13414, n13426, 
        n50_adj_2283, n28_adj_2284, n8_adj_2285, n30_adj_2286, n8_adj_2287, 
        n8_adj_2288, n24212, n24540, n24535, n24532, n24529, n24526, 
        n24523, n24520, n24517, n24514, n24508, n24505, n24502, 
        n24499, n24496, n24493, n24490, n24487, n24469, n24466, 
        n24463, n24460, n24457, n9, n24454, n7, n24431, n24428, 
        n24425, n24422, n49_adj_2289, n24418, n24416, n24413, n24410, 
        n24407, n24404, n24401, n24398, n24394, n24392, n13, n24209, 
        n24203, n24389, n24386, n19, n24367, n24364, n20_adj_2290, 
        n24200, n24197, n24194, n24191, n1_adj_2291, n24350, n24347, 
        n24148, n24188, n23947, n22943, n46_adj_2292, n47_adj_2293, 
        n53_adj_2294, n48_adj_2295, n7584, n24326, n24323, n9513, 
        n8_adj_2296, n24316, n43_adj_2297, n24313, n24310, n44_adj_2298, 
        n24307, n25, n24185, n24182, n24283, n25_adj_2299, n24179;
    
    VCC i2 (.Y(VCC_net));
    lighthouse_ootx_decoder_default ootx_decoder (.\lighthouse[0] (lighthouse[0]), 
            .n6333({Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, 
            Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, 
            n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, 
            Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, 
            Open_19, Open_20, Open_21, Open_22, Open_23}), .counter_from_last_rise({Open_24, 
            Open_25, Open_26, Open_27, Open_28, Open_29, Open_30, 
            Open_31, Open_32, Open_33, Open_34, Open_35, Open_36, 
            counter_from_last_rise[18:13], Open_37, Open_38, Open_39, 
            Open_40, Open_41, Open_42, Open_43, Open_44, counter_from_last_rise[4:0]}), 
            .GND_net(GND_net), .\ootx_payload_o[1][0] (n4568[0]), .clock_c(clock_c), 
            .n1(n1), .n1_adj_1(n1_adj_2267), .n1000(n1000), .data(data), 
            .n1194(n1194), .\ootx_payloads_N_1730[1] (ootx_payloads_N_1730[1]), 
            .n2851({n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
            n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
            n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, 
            n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882}), 
            .bit_counters_0_7(bit_counters_0_7), .bit_counters_1_7(bit_counters_1_7), 
            .bit_counters_0_8(bit_counters_0_8), .bit_counters_1_8(bit_counters_1_8), 
            .bit_counters_0_9(bit_counters_0_9), .bit_counters_1_9(bit_counters_1_9), 
            .\ootx_payloads_N_1730[2] (ootx_payloads_N_1730[2]), .n24018(n24018), 
            .\ootx_payloads_N_1699[4] (ootx_payloads_N_1699[4]), .n13221(n13221), 
            .reset_c(reset_c), .new_data(new_data), .ootx_payloads_N_1744({ootx_payloads_N_1744}), 
            .bit_counters_0_10(bit_counters_0_10), .bit_counters_1_10(bit_counters_1_10), 
            .\ootx_payloads_N_1730[3] (ootx_payloads_N_1730[3]), .n337({n338, 
            n339, n340, n341, n342, n343, n344, n345, n346, 
            n347, n348, n349, n350, n351, n352, n353, n354, 
            n355, n356, n357, n358, n359, n360, n361, n362, 
            n363, n364, n365, n366, n367, n368}), .n998(n998), 
            .n1195(n1195), .n996(n996), .n1196(n1196), .n994(n994), 
            .n1197(n1197), .VCC_net(VCC_net), .n992(n992), .n1198(n1198), 
            .n766(n766), .n1311(n1311), .n13(n13), .n990(n990), .n1199(n1199), 
            .n988(n988), .n1200(n1200), .n1_adj_2(n1_adj_2256), .n9797(n9797), 
            .n23974(n23974), .n8(n8_adj_2280), .bit_counters_0_19(bit_counters_0_19), 
            .bit_counters_1_19(bit_counters_1_19), .n23003(n23003), .data_counters_0_0(data_counters_0_0), 
            .n23005(n23005), .data_counters_0_1(data_counters_0_1), .n23007(n23007), 
            .data_counters_0_2(data_counters_0_2), .n23009(n23009), .data_counters_0_3(data_counters_0_3), 
            .n23011(n23011), .data_counters_0_4(data_counters_0_4), .n23013(n23013), 
            .data_counters_0_5(data_counters_0_5), .n23015(n23015), .data_counters_0_6(data_counters_0_6), 
            .n23017(n23017), .data_counters_0_7(data_counters_0_7), .n23019(n23019), 
            .data_counters_0_8(data_counters_0_8), .n23021(n23021), .data_counters_0_9(data_counters_0_9), 
            .n23023(n23023), .data_counters_0_10(data_counters_0_10), .n1_adj_3(n1_adj_2291), 
            .n23025(n23025), .data_counters_0_11(data_counters_0_11), .n23027(n23027), 
            .data_counters_0_12(data_counters_0_12), .n23029(n23029), .data_counters_0_13(data_counters_0_13), 
            .n23031(n23031), .data_counters_0_14(data_counters_0_14), .n23033(n23033), 
            .data_counters_0_15(data_counters_0_15), .n23035(n23035), .data_counters_0_16(data_counters_0_16), 
            .n23037(n23037), .data_counters_0_17(data_counters_0_17), .n23039(n23039), 
            .data_counters_0_18(data_counters_0_18), .n23041(n23041), .data_counters_0_19(data_counters_0_19), 
            .n23043(n23043), .data_counters_0_20(data_counters_0_20), .n23045(n23045), 
            .data_counters_0_21(data_counters_0_21), .n23047(n23047), .data_counters_0_22(data_counters_0_22), 
            .n23049(n23049), .data_counters_0_23(data_counters_0_23), .n23051(n23051), 
            .data_counters_0_24(data_counters_0_24), .n23053(n23053), .data_counters_0_25(data_counters_0_25), 
            .n23055(n23055), .data_counters_0_26(data_counters_0_26), .n23057(n23057), 
            .data_counters_0_27(data_counters_0_27), .n23059(n23059), .data_counters_0_28(data_counters_0_28), 
            .n23061(n23061), .data_counters_0_29(data_counters_0_29), .n23063(n23063), 
            .data_counters_0_30(data_counters_0_30), .n23065(n23065), .data_counters_1_0(data_counters_1_0), 
            .n23067(n23067), .data_counters_1_1(data_counters_1_1), .n23069(n23069), 
            .data_counters_1_2(data_counters_1_2), .n23071(n23071), .data_counters_1_3(data_counters_1_3), 
            .n23073(n23073), .data_counters_1_4(data_counters_1_4), .n23075(n23075), 
            .data_counters_1_5(data_counters_1_5), .n23077(n23077), .data_counters_1_6(data_counters_1_6), 
            .n23079(n23079), .data_counters_1_7(data_counters_1_7), .n23081(n23081), 
            .data_counters_1_8(data_counters_1_8), .n23083(n23083), .data_counters_1_9(data_counters_1_9), 
            .n23085(n23085), .data_counters_1_10(data_counters_1_10), .n23087(n23087), 
            .data_counters_1_11(data_counters_1_11), .n23089(n23089), .data_counters_1_12(data_counters_1_12), 
            .n23091(n23091), .data_counters_1_13(data_counters_1_13), .n23093(n23093), 
            .data_counters_1_14(data_counters_1_14), .n23095(n23095), .data_counters_1_15(data_counters_1_15), 
            .n23097(n23097), .data_counters_1_16(data_counters_1_16), .n23099(n23099), 
            .data_counters_1_17(data_counters_1_17), .n23101(n23101), .data_counters_1_18(data_counters_1_18), 
            .n23103(n23103), .data_counters_1_19(data_counters_1_19), .n23105(n23105), 
            .data_counters_1_20(data_counters_1_20), .n23107(n23107), .data_counters_1_21(data_counters_1_21), 
            .n23109(n23109), .data_counters_1_22(data_counters_1_22), .n23111(n23111), 
            .data_counters_1_23(data_counters_1_23), .n23113(n23113), .data_counters_1_24(data_counters_1_24), 
            .n23115(n23115), .data_counters_1_25(data_counters_1_25), .n23117(n23117), 
            .data_counters_1_26(data_counters_1_26), .n23119(n23119), .data_counters_1_27(data_counters_1_27), 
            .n23121(n23121), .data_counters_1_28(data_counters_1_28), .n23123(n23123), 
            .data_counters_1_29(data_counters_1_29), .n23125(n23125), .data_counters_1_30(data_counters_1_30), 
            .n23475(n23475), .bit_counters_0_0(bit_counters_0_0), .n23477(n23477), 
            .bit_counters_0_1(bit_counters_0_1), .n23479(n23479), .bit_counters_0_2(bit_counters_0_2), 
            .n23481(n23481), .bit_counters_0_3(bit_counters_0_3), .n23483(n23483), 
            .bit_counters_0_4(bit_counters_0_4), .n23485(n23485), .bit_counters_0_5(bit_counters_0_5), 
            .n23487(n23487), .bit_counters_0_6(bit_counters_0_6), .n23489(n23489), 
            .n23491(n23491), .n23493(n23493), .n23495(n23495), .n23497(n23497), 
            .bit_counters_0_11(bit_counters_0_11), .n23499(n23499), .bit_counters_0_12(bit_counters_0_12), 
            .n23501(n23501), .bit_counters_0_13(bit_counters_0_13), .n23503(n23503), 
            .bit_counters_0_14(bit_counters_0_14), .n23505(n23505), .bit_counters_0_15(bit_counters_0_15), 
            .n23507(n23507), .bit_counters_0_16(bit_counters_0_16), .n23509(n23509), 
            .bit_counters_0_17(bit_counters_0_17), .n23469(n23469), .bit_counters_0_18(bit_counters_0_18), 
            .n23463(n23463), .n23457(n23457), .bit_counters_0_20(bit_counters_0_20), 
            .n23451(n23451), .bit_counters_0_21(bit_counters_0_21), .n23445(n23445), 
            .bit_counters_0_22(bit_counters_0_22), .n23439(n23439), .bit_counters_0_23(bit_counters_0_23), 
            .n23433(n23433), .bit_counters_0_24(bit_counters_0_24), .n23427(n23427), 
            .bit_counters_0_25(bit_counters_0_25), .n23421(n23421), .bit_counters_0_26(bit_counters_0_26), 
            .n23415(n23415), .bit_counters_0_27(bit_counters_0_27), .n23409(n23409), 
            .bit_counters_0_28(bit_counters_0_28), .n23399(n23399), .bit_counters_0_29(bit_counters_0_29), 
            .n23389(n23389), .bit_counters_0_30(bit_counters_0_30), .n23511(n23511), 
            .bit_counters_1_0(bit_counters_1_0), .n23513(n23513), .bit_counters_1_1(bit_counters_1_1), 
            .n23515(n23515), .bit_counters_1_2(bit_counters_1_2), .n23517(n23517), 
            .bit_counters_1_3(bit_counters_1_3), .n23519(n23519), .bit_counters_1_4(bit_counters_1_4), 
            .n23521(n23521), .bit_counters_1_5(bit_counters_1_5), .n23523(n23523), 
            .bit_counters_1_6(bit_counters_1_6), .n23525(n23525), .n23527(n23527), 
            .n23529(n23529), .n23531(n23531), .n23533(n23533), .bit_counters_1_11(bit_counters_1_11), 
            .n23535(n23535), .bit_counters_1_12(bit_counters_1_12), .n23537(n23537), 
            .bit_counters_1_13(bit_counters_1_13), .n23539(n23539), .bit_counters_1_14(bit_counters_1_14), 
            .n23541(n23541), .bit_counters_1_15(bit_counters_1_15), .n23543(n23543), 
            .bit_counters_1_16(bit_counters_1_16), .n23545(n23545), .bit_counters_1_17(bit_counters_1_17), 
            .n23471(n23471), .bit_counters_1_18(bit_counters_1_18), .n23465(n23465), 
            .n23459(n23459), .bit_counters_1_20(bit_counters_1_20), .n23453(n23453), 
            .bit_counters_1_21(bit_counters_1_21), .n23447(n23447), .bit_counters_1_22(bit_counters_1_22), 
            .n23441(n23441), .bit_counters_1_23(bit_counters_1_23), .n23435(n23435), 
            .bit_counters_1_24(bit_counters_1_24), .n23429(n23429), .bit_counters_1_25(bit_counters_1_25), 
            .n23423(n23423), .bit_counters_1_26(bit_counters_1_26), .n23417(n23417), 
            .bit_counters_1_27(bit_counters_1_27), .n986(n986), .n1201(n1201), 
            .n35(n35_adj_2257), .n23411(n23411), .bit_counters_1_28(bit_counters_1_28), 
            .n23401(n23401), .bit_counters_1_29(bit_counters_1_29), .n23391(n23391), 
            .bit_counters_1_30(bit_counters_1_30), .n23697(n23697), .n23639(n23639), 
            .payload_lengths_0_0(payload_lengths_0_0), .n23641(n23641), 
            .payload_lengths_1_0(payload_lengths_1_0), .n8_adj_4(n8_adj_2279), 
            .n8_adj_5(n8_adj_2278), .n8_adj_6(n8_adj_2277), .n2282(n2282), 
            .n8_adj_7(n8_adj_2281), .n984(n984), .n1202(n1202), .n8_adj_8(n8_adj_2296), 
            .\counter_from_last_rise[6] (counter_from_last_rise[6]), .n8_adj_9(n8), 
            .\counter_from_last_rise[7] (counter_from_last_rise[7]), .n8_adj_10(n8_adj_2251), 
            .\counter_from_last_rise[8] (counter_from_last_rise[8]), .n8_adj_11(n8_adj_2265), 
            .\counter_from_last_rise[9] (counter_from_last_rise[9]), .n8_adj_12(n8_adj_2275), 
            .\counter_from_last_rise[10] (counter_from_last_rise[10]), .n8_adj_13(n8_adj_2282), 
            .\counter_from_last_rise[11] (counter_from_last_rise[11]), .n8_adj_14(n8_adj_2285), 
            .\counter_from_last_rise[12] (counter_from_last_rise[12]), .n8_adj_15(n8_adj_2287), 
            .n8_adj_16(n8_adj_2288), .n8_adj_17(n8_adj_2266), .n8_adj_18(n8_adj_2253), 
            .n8_adj_19(n8_adj_2254), .n8_adj_20(n8_adj_2255), .n8_adj_21(n8_adj_2258), 
            .\counter_from_last_rise[19] (counter_from_last_rise[19]), .n8_adj_22(n8_adj_2259), 
            .\counter_from_last_rise[20] (counter_from_last_rise[20]), .n8_adj_23(n8_adj_2260), 
            .\counter_from_last_rise[21] (counter_from_last_rise[21]), .n8_adj_24(n8_adj_2261), 
            .\counter_from_last_rise[22] (counter_from_last_rise[22]), .n8_adj_25(n8_adj_2262), 
            .\counter_from_last_rise[23] (counter_from_last_rise[23]), .n8_adj_26(n8_adj_2263), 
            .\counter_from_last_rise[24] (counter_from_last_rise[24]), .n8_adj_27(n8_adj_2264), 
            .\counter_from_last_rise[25] (counter_from_last_rise[25]), .n8_adj_28(n8_adj_2268), 
            .\counter_from_last_rise[26] (counter_from_last_rise[26]), .n8_adj_29(n8_adj_2269), 
            .\counter_from_last_rise[27] (counter_from_last_rise[27]), .n8_adj_30(n8_adj_2273), 
            .\counter_from_last_rise[28] (counter_from_last_rise[28]), .n8_adj_31(n8_adj_2274), 
            .\counter_from_last_rise[29] (counter_from_last_rise[29]), .n23407(n23407), 
            .\counter_from_last_rise[30] (counter_from_last_rise[30]), .n23397(n23397), 
            .\counter_from_last_rise[31] (counter_from_last_rise[31]), .n12201(n12201), 
            .\ootx_payload_o[0][263] (n4551[263]), .n12200(n12200), .\ootx_payload_o[0][262] (n4551[262]), 
            .n12199(n12199), .\ootx_payload_o[0][261] (n4551[261]), .n12198(n12198), 
            .\ootx_payload_o[0][260] (n4551[260]), .n12197(n12197), .\ootx_payload_o[0][259] (n4551[259]), 
            .n12196(n12196), .\ootx_payload_o[0][258] (n4551[258]), .n12195(n12195), 
            .\ootx_payload_o[0][257] (n4551[257]), .n12194(n12194), .\ootx_payload_o[0][256] (n4551[256]), 
            .n12193(n12193), .\ootx_payload_o[0][255] (n4551[255]), .n12192(n12192), 
            .\ootx_payload_o[0][254] (n4551[254]), .n12191(n12191), .\ootx_payload_o[0][253] (n4551[253]), 
            .n12190(n12190), .\ootx_payload_o[0][252] (n4551[252]), .n12189(n12189), 
            .\ootx_payload_o[0][251] (n4551[251]), .n12188(n12188), .\ootx_payload_o[0][250] (n4551[250]), 
            .n12187(n12187), .\ootx_payload_o[0][249] (n4551[249]), .n12186(n12186), 
            .\ootx_payload_o[0][248] (n4551[248]), .n12185(n12185), .\ootx_payload_o[0][247] (n4551[247]), 
            .n12184(n12184), .\ootx_payload_o[0][246] (n4551[246]), .n12183(n12183), 
            .\ootx_payload_o[0][245] (n4551[245]), .n12182(n12182), .\ootx_payload_o[0][244] (n4551[244]), 
            .n12181(n12181), .\ootx_payload_o[0][243] (n4551[243]), .n12180(n12180), 
            .\ootx_payload_o[0][242] (n4551[242]), .n12179(n12179), .\ootx_payload_o[0][241] (n4551[241]), 
            .n12178(n12178), .\ootx_payload_o[0][240] (n4551[240]), .n12177(n12177), 
            .\ootx_payload_o[0][239] (n4551[239]), .n12176(n12176), .\ootx_payload_o[0][238] (n4551[238]), 
            .n12175(n12175), .\ootx_payload_o[0][237] (n4551[237]), .n12174(n12174), 
            .\ootx_payload_o[0][236] (n4551[236]), .n12173(n12173), .\ootx_payload_o[0][235] (n4551[235]), 
            .n12172(n12172), .\ootx_payload_o[0][234] (n4551[234]), .n12171(n12171), 
            .\ootx_payload_o[0][233] (n4551[233]), .n12170(n12170), .\ootx_payload_o[0][232] (n4551[232]), 
            .n12169(n12169), .\ootx_payload_o[0][231] (n4551[231]), .n12168(n12168), 
            .\ootx_payload_o[0][230] (n4551[230]), .n12167(n12167), .\ootx_payload_o[0][229] (n4551[229]), 
            .n12166(n12166), .\ootx_payload_o[0][228] (n4551[228]), .n12165(n12165), 
            .\ootx_payload_o[0][227] (n4551[227]), .n12164(n12164), .\ootx_payload_o[0][226] (n4551[226]), 
            .n12163(n12163), .\ootx_payload_o[0][225] (n4551[225]), .n12162(n12162), 
            .\ootx_payload_o[0][224] (n4551[224]), .n12161(n12161), .\ootx_payload_o[0][223] (n4551[223]), 
            .n12160(n12160), .\ootx_payload_o[0][222] (n4551[222]), .n12159(n12159), 
            .\ootx_payload_o[0][221] (n4551[221]), .n12158(n12158), .\ootx_payload_o[0][220] (n4551[220]), 
            .n12157(n12157), .\ootx_payload_o[0][219] (n4551[219]), .n12156(n12156), 
            .\ootx_payload_o[0][218] (n4551[218]), .n12155(n12155), .\ootx_payload_o[0][217] (n4551[217]), 
            .n12154(n12154), .\ootx_payload_o[0][216] (n4551[216]), .n12153(n12153), 
            .\ootx_payload_o[0][215] (n4551[215]), .n12152(n12152), .\ootx_payload_o[0][214] (n4551[214]), 
            .n12151(n12151), .\ootx_payload_o[0][213] (n4551[213]), .n12150(n12150), 
            .\ootx_payload_o[0][212] (n4551[212]), .n12149(n12149), .\ootx_payload_o[0][211] (n4551[211]), 
            .n12148(n12148), .\ootx_payload_o[0][210] (n4551[210]), .n12147(n12147), 
            .\ootx_payload_o[0][209] (n4551[209]), .n12146(n12146), .\ootx_payload_o[0][208] (n4551[208]), 
            .n12145(n12145), .\ootx_payload_o[0][207] (n4551[207]), .n12144(n12144), 
            .\ootx_payload_o[0][206] (n4551[206]), .n12143(n12143), .\ootx_payload_o[0][205] (n4551[205]), 
            .n12142(n12142), .\ootx_payload_o[0][204] (n4551[204]), .n12141(n12141), 
            .\ootx_payload_o[0][203] (n4551[203]), .n12140(n12140), .\ootx_payload_o[0][202] (n4551[202]), 
            .n12139(n12139), .\ootx_payload_o[0][201] (n4551[201]), .n12138(n12138), 
            .\ootx_payload_o[0][200] (n4551[200]), .n12137(n12137), .\ootx_payload_o[0][199] (n4551[199]), 
            .n12136(n12136), .\ootx_payload_o[0][198] (n4551[198]), .n12135(n12135), 
            .\ootx_payload_o[0][197] (n4551[197]), .n12134(n12134), .\ootx_payload_o[0][196] (n4551[196]), 
            .n12133(n12133), .\ootx_payload_o[0][195] (n4551[195]), .n12132(n12132), 
            .\ootx_payload_o[0][194] (n4551[194]), .n12131(n12131), .\ootx_payload_o[0][193] (n4551[193]), 
            .n12130(n12130), .\ootx_payload_o[0][192] (n4551[192]), .n12129(n12129), 
            .\ootx_payload_o[0][191] (n4551[191]), .n12128(n12128), .\ootx_payload_o[0][190] (n4551[190]), 
            .n12127(n12127), .\ootx_payload_o[0][189] (n4551[189]), .n12126(n12126), 
            .\ootx_payload_o[0][188] (n4551[188]), .n12125(n12125), .\ootx_payload_o[0][187] (n4551[187]), 
            .n12124(n12124), .\ootx_payload_o[0][186] (n4551[186]), .n12123(n12123), 
            .\ootx_payload_o[0][185] (n4551[185]), .n12122(n12122), .\ootx_payload_o[0][184] (n4551[184]), 
            .n12121(n12121), .\ootx_payload_o[0][183] (n4551[183]), .n12120(n12120), 
            .\ootx_payload_o[0][182] (n4551[182]), .n12119(n12119), .\ootx_payload_o[0][181] (n4551[181]), 
            .n12118(n12118), .\ootx_payload_o[0][180] (n4551[180]), .n12117(n12117), 
            .\ootx_payload_o[0][179] (n4551[179]), .n12116(n12116), .\ootx_payload_o[0][178] (n4551[178]), 
            .n12115(n12115), .\ootx_payload_o[0][177] (n4551[177]), .n12114(n12114), 
            .\ootx_payload_o[0][176] (n4551[176]), .n12113(n12113), .\ootx_payload_o[0][175] (n4551[175]), 
            .n12112(n12112), .\ootx_payload_o[0][174] (n4551[174]), .n12111(n12111), 
            .\ootx_payload_o[0][173] (n4551[173]), .n12110(n12110), .\ootx_payload_o[0][172] (n4551[172]), 
            .n12109(n12109), .\ootx_payload_o[0][171] (n4551[171]), .n12108(n12108), 
            .\ootx_payload_o[0][170] (n4551[170]), .n12107(n12107), .\ootx_payload_o[0][169] (n4551[169]), 
            .n12106(n12106), .\ootx_payload_o[0][168] (n4551[168]), .n12105(n12105), 
            .\ootx_payload_o[0][167] (n4551[167]), .n12104(n12104), .\ootx_payload_o[0][166] (n4551[166]), 
            .n12103(n12103), .\ootx_payload_o[0][165] (n4551[165]), .n12102(n12102), 
            .\ootx_payload_o[0][164] (n4551[164]), .n12101(n12101), .\ootx_payload_o[0][163] (n4551[163]), 
            .n12100(n12100), .\ootx_payload_o[0][162] (n4551[162]), .n12099(n12099), 
            .\ootx_payload_o[0][161] (n4551[161]), .n12098(n12098), .\ootx_payload_o[0][160] (n4551[160]), 
            .n12097(n12097), .\ootx_payload_o[0][159] (n4551[159]), .n12096(n12096), 
            .\ootx_payload_o[0][158] (n4551[158]), .n12095(n12095), .\ootx_payload_o[0][157] (n4551[157]), 
            .n12094(n12094), .\ootx_payload_o[0][156] (n4551[156]), .n12093(n12093), 
            .\ootx_payload_o[0][155] (n4551[155]), .n12092(n12092), .\ootx_payload_o[0][154] (n4551[154]), 
            .n12091(n12091), .\ootx_payload_o[0][153] (n4551[153]), .n12090(n12090), 
            .\ootx_payload_o[0][152] (n4551[152]), .n12089(n12089), .\ootx_payload_o[0][151] (n4551[151]), 
            .n12088(n12088), .\ootx_payload_o[0][150] (n4551[150]), .n12087(n12087), 
            .\ootx_payload_o[0][149] (n4551[149]), .n12086(n12086), .\ootx_payload_o[0][148] (n4551[148]), 
            .n12085(n12085), .\ootx_payload_o[0][147] (n4551[147]), .n12084(n12084), 
            .\ootx_payload_o[0][146] (n4551[146]), .n12083(n12083), .\ootx_payload_o[0][145] (n4551[145]), 
            .n12082(n12082), .\ootx_payload_o[0][144] (n4551[144]), .n12081(n12081), 
            .\ootx_payload_o[0][143] (n4551[143]), .n12080(n12080), .\ootx_payload_o[0][142] (n4551[142]), 
            .n12079(n12079), .\ootx_payload_o[0][141] (n4551[141]), .n12078(n12078), 
            .\ootx_payload_o[0][140] (n4551[140]), .n12077(n12077), .\ootx_payload_o[0][139] (n4551[139]), 
            .n12076(n12076), .\ootx_payload_o[0][138] (n4551[138]), .n12075(n12075), 
            .\ootx_payload_o[0][137] (n4551[137]), .n12074(n12074), .\ootx_payload_o[0][136] (n4551[136]), 
            .n12073(n12073), .\ootx_payload_o[0][135] (n4551[135]), .n12072(n12072), 
            .\ootx_payload_o[0][134] (n4551[134]), .n12071(n12071), .\ootx_payload_o[0][133] (n4551[133]), 
            .n12070(n12070), .\ootx_payload_o[0][132] (n4551[132]), .n12069(n12069), 
            .\ootx_payload_o[0][131] (n4551[131]), .n12068(n12068), .\ootx_payload_o[0][130] (n4551[130]), 
            .n12067(n12067), .\ootx_payload_o[0][129] (n4551[129]), .n12066(n12066), 
            .\ootx_payload_o[0][128] (n4551[128]), .n12065(n12065), .\ootx_payload_o[0][127] (n4551[127]), 
            .n12064(n12064), .\ootx_payload_o[0][126] (n4551[126]), .n12063(n12063), 
            .\ootx_payload_o[0][125] (n4551[125]), .n12062(n12062), .\ootx_payload_o[0][124] (n4551[124]), 
            .n12061(n12061), .\ootx_payload_o[0][123] (n4551[123]), .n12060(n12060), 
            .\ootx_payload_o[0][122] (n4551[122]), .n12059(n12059), .\ootx_payload_o[0][121] (n4551[121]), 
            .n12058(n12058), .\ootx_payload_o[0][120] (n4551[120]), .n12057(n12057), 
            .\ootx_payload_o[0][119] (n4551[119]), .n12056(n12056), .\ootx_payload_o[0][118] (n4551[118]), 
            .n12055(n12055), .\ootx_payload_o[0][117] (n4551[117]), .n12054(n12054), 
            .\ootx_payload_o[0][116] (n4551[116]), .n12053(n12053), .\ootx_payload_o[0][115] (n4551[115]), 
            .n12052(n12052), .\ootx_payload_o[0][114] (n4551[114]), .n12051(n12051), 
            .\ootx_payload_o[0][113] (n4551[113]), .n12050(n12050), .\ootx_payload_o[0][112] (n4551[112]), 
            .n12049(n12049), .\ootx_payload_o[0][111] (n4551[111]), .n12048(n12048), 
            .\ootx_payload_o[0][110] (n4551[110]), .n12047(n12047), .\ootx_payload_o[0][109] (n4551[109]), 
            .n12046(n12046), .\ootx_payload_o[0][108] (n4551[108]), .n12045(n12045), 
            .\ootx_payload_o[0][107] (n4551[107]), .n12044(n12044), .\ootx_payload_o[0][106] (n4551[106]), 
            .n12043(n12043), .\ootx_payload_o[0][105] (n4551[105]), .n12042(n12042), 
            .\ootx_payload_o[0][104] (n4551[104]), .n12041(n12041), .\ootx_payload_o[0][103] (n4551[103]), 
            .n12040(n12040), .\ootx_payload_o[0][102] (n4551[102]), .n12039(n12039), 
            .\ootx_payload_o[0][101] (n4551[101]), .n12038(n12038), .\ootx_payload_o[0][100] (n4551[100]), 
            .n12037(n12037), .\ootx_payload_o[0][99] (n4551[99]), .n12036(n12036), 
            .\ootx_payload_o[0][98] (n4551[98]), .n12035(n12035), .\ootx_payload_o[0][97] (n4551[97]), 
            .n12034(n12034), .\ootx_payload_o[0][96] (n4551[96]), .n12033(n12033), 
            .\ootx_payload_o[0][95] (n4551[95]), .n12032(n12032), .\ootx_payload_o[0][94] (n4551[94]), 
            .n12031(n12031), .\ootx_payload_o[0][93] (n4551[93]), .n12030(n12030), 
            .\ootx_payload_o[0][92] (n4551[92]), .n12029(n12029), .\ootx_payload_o[0][91] (n4551[91]), 
            .n12028(n12028), .\ootx_payload_o[0][90] (n4551[90]), .n12027(n12027), 
            .\ootx_payload_o[0][89] (n4551[89]), .n12026(n12026), .\ootx_payload_o[0][88] (n4551[88]), 
            .n12025(n12025), .\ootx_payload_o[0][87] (n4551[87]), .n12024(n12024), 
            .\ootx_payload_o[0][86] (n4551[86]), .n12023(n12023), .\ootx_payload_o[0][85] (n4551[85]), 
            .n12022(n12022), .\ootx_payload_o[0][84] (n4551[84]), .n12021(n12021), 
            .\ootx_payload_o[0][83] (n4551[83]), .n12020(n12020), .\ootx_payload_o[0][82] (n4551[82]), 
            .n12019(n12019), .\ootx_payload_o[0][81] (n4551[81]), .n12018(n12018), 
            .\ootx_payload_o[0][80] (n4551[80]), .n12017(n12017), .\ootx_payload_o[0][79] (n4551[79]), 
            .n12016(n12016), .\ootx_payload_o[0][78] (n4551[78]), .n12015(n12015), 
            .\ootx_payload_o[0][77] (n4551[77]), .n12014(n12014), .\ootx_payload_o[0][76] (n4551[76]), 
            .n12013(n12013), .\ootx_payload_o[0][75] (n4551[75]), .n12012(n12012), 
            .\ootx_payload_o[0][74] (n4551[74]), .n12011(n12011), .\ootx_payload_o[0][73] (n4551[73]), 
            .n12010(n12010), .\ootx_payload_o[0][72] (n4551[72]), .n12009(n12009), 
            .\ootx_payload_o[0][71] (n4551[71]), .n12008(n12008), .\ootx_payload_o[0][70] (n4551[70]), 
            .n12007(n12007), .\ootx_payload_o[0][69] (n4551[69]), .n12006(n12006), 
            .\ootx_payload_o[0][68] (n4551[68]), .n12005(n12005), .\ootx_payload_o[0][67] (n4551[67]), 
            .n12004(n12004), .\ootx_payload_o[0][66] (n4551[66]), .n12003(n12003), 
            .\ootx_payload_o[0][65] (n4551[65]), .n12002(n12002), .\ootx_payload_o[0][64] (n4551[64]), 
            .n12001(n12001), .\ootx_payload_o[0][63] (n4551[63]), .n12000(n12000), 
            .\ootx_payload_o[0][62] (n4551[62]), .n11999(n11999), .\ootx_payload_o[0][61] (n4551[61]), 
            .n11998(n11998), .\ootx_payload_o[0][60] (n4551[60]), .n11997(n11997), 
            .\ootx_payload_o[0][59] (n4551[59]), .n11996(n11996), .\ootx_payload_o[0][58] (n4551[58]), 
            .n11995(n11995), .\ootx_payload_o[0][57] (n4551[57]), .n11994(n11994), 
            .\ootx_payload_o[0][56] (n4551[56]), .n11993(n11993), .\ootx_payload_o[0][55] (n4551[55]), 
            .n11992(n11992), .\ootx_payload_o[0][54] (n4551[54]), .n11991(n11991), 
            .\ootx_payload_o[0][53] (n4551[53]), .n11990(n11990), .\ootx_payload_o[0][52] (n4551[52]), 
            .n938(n938), .n1225(n1225), .n11989(n11989), .\ootx_payload_o[0][51] (n4551[51]), 
            .n11988(n11988), .\ootx_payload_o[0][50] (n4551[50]), .n11987(n11987), 
            .\ootx_payload_o[0][49] (n4551[49]), .n11986(n11986), .\ootx_payload_o[0][48] (n4551[48]), 
            .n11985(n11985), .\ootx_payload_o[0][47] (n4551[47]), .n11984(n11984), 
            .\ootx_payload_o[0][46] (n4551[46]), .n11983(n11983), .\ootx_payload_o[0][45] (n4551[45]), 
            .n958(n958), .n1215(n1215), .n11982(n11982), .\ootx_payload_o[0][44] (n4551[44]), 
            .n30(n30_adj_2286), .n11981(n11981), .\ootx_payload_o[0][43] (n4551[43]), 
            .n11980(n11980), .\ootx_payload_o[0][42] (n4551[42]), .n11979(n11979), 
            .\ootx_payload_o[0][41] (n4551[41]), .n11978(n11978), .\ootx_payload_o[0][40] (n4551[40]), 
            .n11977(n11977), .\ootx_payload_o[0][39] (n4551[39]), .n982(n982), 
            .n1203(n1203), .n11976(n11976), .\ootx_payload_o[0][38] (n4551[38]), 
            .n11975(n11975), .\ootx_payload_o[0][37] (n4551[37]), .n11974(n11974), 
            .\ootx_payload_o[0][36] (n4551[36]), .n11973(n11973), .\ootx_payload_o[0][35] (n4551[35]), 
            .sensor_state(sensor_state), .n11972(n11972), .\ootx_payload_o[0][34] (n4551[34]), 
            .n11971(n11971), .\ootx_payload_o[0][33] (n4551[33]), .n11970(n11970), 
            .\ootx_payload_o[0][32] (n4551[32]), .n11969(n11969), .\ootx_payload_o[0][31] (n4551[31]), 
            .n11968(n11968), .\ootx_payload_o[0][30] (n4551[30]), .n11967(n11967), 
            .\ootx_payload_o[0][29] (n4551[29]), .n11966(n11966), .\ootx_payload_o[0][28] (n4551[28]), 
            .n11965(n11965), .\ootx_payload_o[0][27] (n4551[27]), .n11964(n11964), 
            .\ootx_payload_o[0][26] (n4551[26]), .n11963(n11963), .\ootx_payload_o[0][25] (n4551[25]), 
            .n11962(n11962), .\ootx_payload_o[0][24] (n4551[24]), .n11961(n11961), 
            .\ootx_payload_o[0][23] (n4551[23]), .n11960(n11960), .\ootx_payload_o[0][22] (n4551[22]), 
            .n11959(n11959), .\ootx_payload_o[0][21] (n4551[21]), .n680(n680), 
            .n1354(n1354), .n712(n712), .n1338(n1338), .\ootx_payloads_N_1699[5] (ootx_payloads_N_1699[5]), 
            .\ootx_payloads_N_1699[3] (ootx_payloads_N_1699[3]), .\ootx_payloads_N_1699[15] (ootx_payloads_N_1699[15]), 
            .n34({n35, n36}), .n11958(n11958), .\ootx_payload_o[0][20] (n4551[20]), 
            .n11957(n11957), .\ootx_payload_o[0][19] (n4551[19]), .n11956(n11956), 
            .\ootx_payload_o[0][18] (n4551[18]), .n11955(n11955), .\ootx_payload_o[0][17] (n4551[17]), 
            .n11954(n11954), .\ootx_payload_o[0][16] (n4551[16]), .n11953(n11953), 
            .\ootx_payload_o[0][15] (n4551[15]), .n11952(n11952), .\ootx_payload_o[0][14] (n4551[14]), 
            .n11951(n11951), .\ootx_payload_o[0][13] (n4551[13]), .n11950(n11950), 
            .\ootx_payload_o[0][12] (n4551[12]), .n11949(n11949), .\ootx_payload_o[0][11] (n4551[11]), 
            .n11948(n11948), .\ootx_payload_o[0][10] (n4551[10]), .n11947(n11947), 
            .\ootx_payload_o[0][9] (n4551[9]), .n11946(n11946), .\ootx_payload_o[0][8] (n4551[8]), 
            .n11945(n11945), .\ootx_payload_o[0][7] (n4551[7]), .n11944(n11944), 
            .\ootx_payload_o[0][6] (n4551[6]), .n11943(n11943), .\ootx_payload_o[0][5] (n4551[5]), 
            .n11942(n11942), .\ootx_payload_o[0][4] (n4551[4]), .n11941(n11941), 
            .\ootx_payload_o[0][3] (n4551[3]), .n11940(n11940), .\ootx_payload_o[0][2] (n4551[2]), 
            .n11939(n11939), .\ootx_payload_o[0][1] (n4551[1]), .\ootx_crc32_o[1] ({\ootx_crc32_o[1] }), 
            .\ootx_crc32_o[0] ({\ootx_crc32_o[0] }), .n1170(n1170), .n1171(n1171), 
            .n1172(n1172), .n1173(n1173), .n1174(n1174), .n1175(n1175), 
            .n1176(n1176), .n1177(n1177), .n1178(n1178), .n1179(n1179), 
            .n1180(n1180), .n1181(n1181), .n1182(n1182), .n1183(n1183), 
            .n1184(n1184), .n1185(n1185), .n1186(n1186), .n1187(n1187), 
            .n1188(n1188), .n1189(n1189), .n1190(n1190), .n1191(n1191), 
            .n1192(n1192), .n1193(n1193), .n640(n640), .n1374(n1374), 
            .n724(n724), .n928(n928), .n1230(n1230), .n1204(n1204), 
            .n1205(n1205), .n1206(n1206), .n1207(n1207), .n1208(n1208), 
            .n1209(n1209), .n1210(n1210), .n1332(n1332), .n1211(n1211), 
            .n1212(n1212), .n1213(n1213), .\ootx_payloads_N_1699[6] (ootx_payloads_N_1699[6]), 
            .\ootx_payloads_N_1699[7] (ootx_payloads_N_1699[7]), .\ootx_payloads_N_1699[8] (ootx_payloads_N_1699[8]), 
            .n1010(n1010), .n1214(n1214), .n754(n754), .n764(n764), 
            .n672(n672), .\ootx_states[0] ({\ootx_states[0] }), .n638(n638), 
            .n1375(n1375), .ootx_payloads_1_263(ootx_payloads_1_263), .n926(n926), 
            .n1231(n1231), .n670(n670), .n1312(n1312), .n20(n20_adj_2290), 
            .ootx_payloads_1_262(ootx_payloads_1_262), .n924(n924), .n1232(n1232), 
            .n636(n636), .n1376(n1376), .n668(n668), .n922(n922), .n1233(n1233), 
            .n634(n634), .n1377(n1377), .n666(n666), .n920(n920), .n1234(n1234), 
            .n632(n632), .n1378(n1378), .n664(n664), .n918(n918), .n1235(n1235), 
            .n662(n662), .n916(n916), .n1236(n1236), .n752(n752), .n1318(n1318), 
            .n660(n660), .n914(n914), .n1237(n1237), .n658(n658), .n678(n678), 
            .n1355(n1355), .n912(n912), .n1238(n1238), .n630(n630), 
            .n1379(n1379), .ootx_payloads_1_261(ootx_payloads_1_261), .ootx_payloads_1_260(ootx_payloads_1_260), 
            .n656(n656), .ootx_payloads_1_259(ootx_payloads_1_259), .n910(n910), 
            .n1239(n1239), .n654(n654), .n1008(n1008), .n676(n676), 
            .n1356(n1356), .n908(n908), .n1240(n1240), .ootx_payloads_1_258(ootx_payloads_1_258), 
            .ootx_payloads_1_257(ootx_payloads_1_257), .ootx_payloads_1_256(ootx_payloads_1_256), 
            .n628(n628), .n1380(n1380), .ootx_payloads_1_255(ootx_payloads_1_255), 
            .\ootx_payloads_N_1699[30] (ootx_payloads_N_1699[30]), .n9200(n9200), 
            .\ootx_payloads_N_1699[9] (ootx_payloads_N_1699[9]), .\ootx_payloads_N_1699[13] (ootx_payloads_N_1699[13]), 
            .\ootx_payloads_N_1699[12] (ootx_payloads_N_1699[12]), .\ootx_payloads_N_1699[11] (ootx_payloads_N_1699[11]), 
            .ootx_payloads_1_254(ootx_payloads_1_254), .ootx_payloads_1_253(ootx_payloads_1_253), 
            .ootx_payloads_1_252(ootx_payloads_1_252), .ootx_payloads_1_251(ootx_payloads_1_251), 
            .n652(n652), .n906(n906), .n1241(n1241), .ootx_payloads_1_250(ootx_payloads_1_250), 
            .ootx_payloads_1_249(ootx_payloads_1_249), .\ootx_payloads_N_1699[10] (ootx_payloads_N_1699[10]), 
            .\ootx_payloads_N_1699[14] (ootx_payloads_N_1699[14]), .n650(n650), 
            .n626(n626), .n1381(n1381), .n904(n904), .n1242(n1242), 
            .n648(n648), .n980(n980), .n624(n624), .n1382(n1382), .ootx_payloads_1_248(ootx_payloads_1_248), 
            .ootx_payloads_1_247(ootx_payloads_1_247), .n902(n902), .n1243(n1243), 
            .n900(n900), .n1244(n1244), .n978(n978), .n674(n674), .n1357(n1357), 
            .n19(n19), .n622(n622), .n1383(n1383), .ootx_payloads_1_246(ootx_payloads_1_246), 
            .ootx_payloads_1_245(ootx_payloads_1_245), .n898(n898), .n1245(n1245), 
            .ootx_payloads_1_244(ootx_payloads_1_244), .n896(n896), .n1246(n1246), 
            .n620(n620), .n1384(n1384), .n6355(n6355), .n894(n894), 
            .n1247(n1247), .n6356(n6356), .n6357(n6357), .\ootx_payloads_N_1730[4] (ootx_payloads_N_1730[4]), 
            .n6358(n6358), .n750(n750), .n1319(n1319), .n618(n618), 
            .n1385(n1385), .n892(n892), .n1248(n1248), .n6359(n6359), 
            .ootx_payloads_1_243(ootx_payloads_1_243), .n6361(n6361), .n890(n890), 
            .n1249(n1249), .ootx_payloads_1_242(ootx_payloads_1_242), .n6362(n6362), 
            .n616(n616), .n1386(n1386), .ootx_payloads_1_241(ootx_payloads_1_241), 
            .ootx_payloads_1_240(ootx_payloads_1_240), .ootx_payloads_1_239(ootx_payloads_1_239), 
            .n1006(n1006), .n888(n888), .n1250(n1250), .ootx_payloads_1_238(ootx_payloads_1_238), 
            .ootx_payloads_1_237(ootx_payloads_1_237), .n886(n886), .n1251(n1251), 
            .n614(n614), .n1387(n1387), .n22943(n22943), .n976(n976), 
            .ootx_payloads_1_236(ootx_payloads_1_236), .n884(n884), .n1252(n1252), 
            .ootx_payloads_1_235(ootx_payloads_1_235), .n882(n882), .n1253(n1253), 
            .ootx_payloads_1_234(ootx_payloads_1_234), .n1358(n1358), .n612(n612), 
            .n1388(n1388), .n880(n880), .n1254(n1254), .n748(n748), 
            .n1320(n1320), .n974(n974), .n878(n878), .n1255(n1255), 
            .n1004(n1004), .n13329(n13329), .data_N_1808(data_N_1808), 
            .n6363(n6363), .n6364(n6364), .n6365(n6365), .ootx_payloads_1_233(ootx_payloads_1_233), 
            .sensor_N_132(sensor_N_132), .n876(n876), .n1256(n1256), .ootx_payloads_1_232(ootx_payloads_1_232), 
            .n610(n610), .n1389(n1389), .ootx_payloads_1_231(ootx_payloads_1_231), 
            .n874(n874), .n1257(n1257), .n872(n872), .n1258(n1258), 
            .n608(n608), .n1390(n1390), .n870(n870), .n1259(n1259), 
            .n746(n746), .n1321(n1321), .n606(n606), .n1391(n1391), 
            .n604(n604), .n1392(n1392), .n710(n710), .n1339(n1339), 
            .n966(n966), .n868(n868), .n1260(n1260), .n602(n602), .n1393(n1393), 
            .n744(n744), .n1322(n1322), .n866(n866), .n1261(n1261), 
            .n600(n600), .n1394(n1394), .n864(n864), .n1262(n1262), 
            .n598(n598), .n1395(n1395), .ootx_payloads_1_230(ootx_payloads_1_230), 
            .ootx_payloads_1_229(ootx_payloads_1_229), .ootx_payloads_1_228(ootx_payloads_1_228), 
            .ootx_payloads_1_227(ootx_payloads_1_227), .n596(n596), .n1396(n1396), 
            .n594(n594), .n1397(n1397), .ootx_payloads_1_226(ootx_payloads_1_226), 
            .ootx_payloads_1_225(ootx_payloads_1_225), .ootx_payloads_1_224(ootx_payloads_1_224), 
            .n592(n592), .n1398(n1398), .ootx_payloads_1_223(ootx_payloads_1_223), 
            .n742(n742), .n1323(n1323), .n862(n862), .n1263(n1263), 
            .n590(n590), .n1399(n1399), .ootx_payloads_1_222(ootx_payloads_1_222), 
            .ootx_payloads_1_221(ootx_payloads_1_221), .\ootx_payload_o[1][1] (n4568[1]), 
            .ootx_payloads_1_220(ootx_payloads_1_220), .ootx_payloads_1_219(ootx_payloads_1_219), 
            .ootx_payloads_1_218(ootx_payloads_1_218), .n588(n588), .n1400(n1400), 
            .ootx_payloads_1_217(ootx_payloads_1_217), .ootx_payloads_1_216(ootx_payloads_1_216), 
            .\ootx_payload_o[1][2] (n4568[2]), .\ootx_payload_o[1][3] (n4568[3]), 
            .\ootx_payload_o[1][4] (n4568[4]), .\ootx_payload_o[1][5] (n4568[5]), 
            .\ootx_payload_o[1][6] (n4568[6]), .\ootx_payload_o[1][7] (n4568[7]), 
            .\ootx_payload_o[1][8] (n4568[8]), .\ootx_payload_o[1][9] (n4568[9]), 
            .\ootx_payload_o[1][10] (n4568[10]), .\ootx_payload_o[1][11] (n4568[11]), 
            .\ootx_payload_o[1][12] (n4568[12]), .\ootx_payload_o[1][13] (n4568[13]), 
            .\ootx_payload_o[1][14] (n4568[14]), .\ootx_payload_o[1][15] (n4568[15]), 
            .\ootx_payload_o[1][16] (n4568[16]), .\ootx_payload_o[1][17] (n4568[17]), 
            .\ootx_payload_o[1][18] (n4568[18]), .\ootx_payload_o[1][19] (n4568[19]), 
            .\ootx_payload_o[1][20] (n4568[20]), .\ootx_payload_o[1][21] (n4568[21]), 
            .\ootx_payload_o[1][22] (n4568[22]), .\ootx_payload_o[1][23] (n4568[23]), 
            .\ootx_payload_o[1][24] (n4568[24]), .\ootx_payload_o[1][25] (n4568[25]), 
            .\ootx_payload_o[1][26] (n4568[26]), .\ootx_payload_o[1][27] (n4568[27]), 
            .\ootx_payload_o[1][28] (n4568[28]), .\ootx_payload_o[1][29] (n4568[29]), 
            .\ootx_payload_o[1][30] (n4568[30]), .\ootx_payload_o[1][31] (n4568[31]), 
            .\ootx_payload_o[1][32] (n4568[32]), .\ootx_payload_o[1][33] (n4568[33]), 
            .\ootx_payload_o[1][34] (n4568[34]), .\ootx_payload_o[1][35] (n4568[35]), 
            .\ootx_payload_o[1][36] (n4568[36]), .\ootx_payload_o[1][37] (n4568[37]), 
            .\ootx_payload_o[1][38] (n4568[38]), .\ootx_payload_o[1][39] (n4568[39]), 
            .\ootx_payload_o[1][40] (n4568[40]), .\ootx_payload_o[1][41] (n4568[41]), 
            .\ootx_payload_o[1][42] (n4568[42]), .\ootx_payload_o[1][43] (n4568[43]), 
            .\ootx_payload_o[1][44] (n4568[44]), .\ootx_payload_o[1][45] (n4568[45]), 
            .\ootx_payload_o[1][46] (n4568[46]), .\ootx_payload_o[1][47] (n4568[47]), 
            .\ootx_payload_o[1][48] (n4568[48]), .\ootx_payload_o[1][49] (n4568[49]), 
            .\ootx_payload_o[1][50] (n4568[50]), .\ootx_payload_o[1][51] (n4568[51]), 
            .\ootx_payload_o[1][52] (n4568[52]), .\ootx_payload_o[1][53] (n4568[53]), 
            .\ootx_payload_o[1][54] (n4568[54]), .\ootx_payload_o[1][55] (n4568[55]), 
            .\ootx_payload_o[1][56] (n4568[56]), .\ootx_payload_o[1][57] (n4568[57]), 
            .\ootx_payload_o[1][58] (n4568[58]), .\ootx_payload_o[1][59] (n4568[59]), 
            .\ootx_payload_o[1][60] (n4568[60]), .\ootx_payload_o[1][61] (n4568[61]), 
            .\ootx_payload_o[1][62] (n4568[62]), .\ootx_payload_o[1][63] (n4568[63]), 
            .\ootx_payload_o[1][64] (n4568[64]), .\ootx_payload_o[1][65] (n4568[65]), 
            .\ootx_payload_o[1][66] (n4568[66]), .\ootx_payload_o[1][67] (n4568[67]), 
            .\ootx_payload_o[1][68] (n4568[68]), .\ootx_payload_o[1][69] (n4568[69]), 
            .\ootx_payload_o[1][70] (n4568[70]), .\ootx_payload_o[1][71] (n4568[71]), 
            .\ootx_payload_o[1][72] (n4568[72]), .\ootx_payload_o[1][73] (n4568[73]), 
            .\ootx_payload_o[1][74] (n4568[74]), .\ootx_payload_o[1][75] (n4568[75]), 
            .\ootx_payload_o[1][76] (n4568[76]), .\ootx_payload_o[1][77] (n4568[77]), 
            .\ootx_payload_o[1][78] (n4568[78]), .\ootx_payload_o[1][79] (n4568[79]), 
            .\ootx_payload_o[1][80] (n4568[80]), .\ootx_payload_o[1][81] (n4568[81]), 
            .\ootx_payload_o[1][82] (n4568[82]), .\ootx_payload_o[1][83] (n4568[83]), 
            .\ootx_payload_o[1][84] (n4568[84]), .\ootx_payload_o[1][85] (n4568[85]), 
            .\ootx_payload_o[1][86] (n4568[86]), .\ootx_payload_o[1][87] (n4568[87]), 
            .\ootx_payload_o[1][88] (n4568[88]), .\ootx_payload_o[1][89] (n4568[89]), 
            .\ootx_payload_o[1][90] (n4568[90]), .\ootx_payload_o[1][91] (n4568[91]), 
            .\ootx_payload_o[1][92] (n4568[92]), .\ootx_payload_o[1][93] (n4568[93]), 
            .\ootx_payload_o[1][94] (n4568[94]), .\ootx_payload_o[1][95] (n4568[95]), 
            .\ootx_payload_o[1][96] (n4568[96]), .\ootx_payload_o[1][97] (n4568[97]), 
            .\ootx_payload_o[1][98] (n4568[98]), .\ootx_payload_o[1][99] (n4568[99]), 
            .\ootx_payload_o[1][100] (n4568[100]), .\ootx_payload_o[1][101] (n4568[101]), 
            .\ootx_payload_o[1][102] (n4568[102]), .\ootx_payload_o[1][103] (n4568[103]), 
            .\ootx_payload_o[1][104] (n4568[104]), .\ootx_payload_o[1][105] (n4568[105]), 
            .\ootx_payload_o[1][106] (n4568[106]), .\ootx_payload_o[1][107] (n4568[107]), 
            .\ootx_payload_o[1][108] (n4568[108]), .\ootx_payload_o[1][109] (n4568[109]), 
            .\ootx_payload_o[1][110] (n4568[110]), .\ootx_payload_o[1][111] (n4568[111]), 
            .\ootx_payload_o[1][112] (n4568[112]), .\ootx_payload_o[1][113] (n4568[113]), 
            .\ootx_payload_o[1][114] (n4568[114]), .\ootx_payload_o[1][115] (n4568[115]), 
            .\ootx_payload_o[1][116] (n4568[116]), .\ootx_payload_o[1][117] (n4568[117]), 
            .\ootx_payload_o[1][118] (n4568[118]), .\ootx_payload_o[1][119] (n4568[119]), 
            .\ootx_payload_o[1][120] (n4568[120]), .\ootx_payload_o[1][121] (n4568[121]), 
            .\ootx_payload_o[1][122] (n4568[122]), .\ootx_payload_o[1][123] (n4568[123]), 
            .\ootx_payload_o[1][124] (n4568[124]), .\ootx_payload_o[1][125] (n4568[125]), 
            .\ootx_payload_o[1][126] (n4568[126]), .\ootx_payload_o[1][127] (n4568[127]), 
            .\ootx_payload_o[1][128] (n4568[128]), .\ootx_payload_o[1][129] (n4568[129]), 
            .\ootx_payload_o[1][130] (n4568[130]), .\ootx_payload_o[1][131] (n4568[131]), 
            .\ootx_payload_o[1][132] (n4568[132]), .\ootx_payload_o[1][133] (n4568[133]), 
            .\ootx_payload_o[1][134] (n4568[134]), .\ootx_payload_o[1][135] (n4568[135]), 
            .\ootx_payload_o[1][136] (n4568[136]), .\ootx_payload_o[1][137] (n4568[137]), 
            .\ootx_payload_o[1][138] (n4568[138]), .\ootx_payload_o[1][139] (n4568[139]), 
            .\ootx_payload_o[1][140] (n4568[140]), .\ootx_payload_o[1][141] (n4568[141]), 
            .\ootx_payload_o[1][142] (n4568[142]), .\ootx_payload_o[1][143] (n4568[143]), 
            .\ootx_payload_o[1][144] (n4568[144]), .\ootx_payload_o[1][145] (n4568[145]), 
            .\ootx_payload_o[1][146] (n4568[146]), .\ootx_payload_o[1][147] (n4568[147]), 
            .\ootx_payload_o[1][148] (n4568[148]), .\ootx_payload_o[1][149] (n4568[149]), 
            .\ootx_payload_o[1][150] (n4568[150]), .\ootx_payload_o[1][151] (n4568[151]), 
            .\ootx_payload_o[1][152] (n4568[152]), .\ootx_payload_o[1][153] (n4568[153]), 
            .\ootx_payload_o[1][154] (n4568[154]), .\ootx_payload_o[1][155] (n4568[155]), 
            .\ootx_payload_o[1][156] (n4568[156]), .\ootx_payload_o[1][157] (n4568[157]), 
            .\ootx_payload_o[1][158] (n4568[158]), .\ootx_payload_o[1][159] (n4568[159]), 
            .\ootx_payload_o[1][160] (n4568[160]), .\ootx_payload_o[1][161] (n4568[161]), 
            .\ootx_payload_o[1][162] (n4568[162]), .\ootx_payload_o[1][163] (n4568[163]), 
            .\ootx_payload_o[1][164] (n4568[164]), .\ootx_payload_o[1][165] (n4568[165]), 
            .\ootx_payload_o[1][166] (n4568[166]), .\ootx_payload_o[1][167] (n4568[167]), 
            .\ootx_payload_o[1][168] (n4568[168]), .\ootx_payload_o[1][169] (n4568[169]), 
            .\ootx_payload_o[1][170] (n4568[170]), .\ootx_payload_o[1][171] (n4568[171]), 
            .\ootx_payload_o[1][172] (n4568[172]), .\ootx_payload_o[1][173] (n4568[173]), 
            .\ootx_payload_o[1][174] (n4568[174]), .\ootx_payload_o[1][175] (n4568[175]), 
            .\ootx_payload_o[1][176] (n4568[176]), .\ootx_payload_o[1][177] (n4568[177]), 
            .\ootx_payload_o[1][178] (n4568[178]), .\ootx_payload_o[1][179] (n4568[179]), 
            .\ootx_payload_o[1][180] (n4568[180]), .\ootx_payload_o[1][181] (n4568[181]), 
            .\ootx_payload_o[1][182] (n4568[182]), .\ootx_payload_o[1][183] (n4568[183]), 
            .\ootx_payload_o[1][184] (n4568[184]), .\ootx_payload_o[1][185] (n4568[185]), 
            .\ootx_payload_o[1][186] (n4568[186]), .\ootx_payload_o[1][187] (n4568[187]), 
            .\ootx_payload_o[1][188] (n4568[188]), .\ootx_payload_o[1][189] (n4568[189]), 
            .\ootx_payload_o[1][190] (n4568[190]), .\ootx_payload_o[1][191] (n4568[191]), 
            .\ootx_payload_o[1][192] (n4568[192]), .\ootx_payload_o[1][193] (n4568[193]), 
            .\ootx_payload_o[1][194] (n4568[194]), .\ootx_payload_o[1][195] (n4568[195]), 
            .\ootx_payload_o[1][196] (n4568[196]), .\ootx_payload_o[1][197] (n4568[197]), 
            .\ootx_payload_o[1][198] (n4568[198]), .\ootx_payload_o[1][199] (n4568[199]), 
            .\ootx_payload_o[1][200] (n4568[200]), .\ootx_payload_o[1][201] (n4568[201]), 
            .\ootx_payload_o[1][202] (n4568[202]), .\ootx_payload_o[1][203] (n4568[203]), 
            .\ootx_payload_o[1][204] (n4568[204]), .\ootx_payload_o[1][205] (n4568[205]), 
            .\ootx_payload_o[1][206] (n4568[206]), .\ootx_payload_o[1][207] (n4568[207]), 
            .\ootx_payload_o[1][208] (n4568[208]), .\ootx_payload_o[1][209] (n4568[209]), 
            .\ootx_payload_o[1][210] (n4568[210]), .\ootx_payload_o[1][211] (n4568[211]), 
            .\ootx_payload_o[1][212] (n4568[212]), .\ootx_payload_o[1][213] (n4568[213]), 
            .\ootx_payload_o[1][214] (n4568[214]), .\ootx_payload_o[1][215] (n4568[215]), 
            .\ootx_payload_o[1][216] (n4568[216]), .\ootx_payload_o[1][217] (n4568[217]), 
            .\ootx_payload_o[1][218] (n4568[218]), .\ootx_payload_o[1][219] (n4568[219]), 
            .\ootx_payload_o[1][220] (n4568[220]), .\ootx_payload_o[1][221] (n4568[221]), 
            .\ootx_payload_o[1][222] (n4568[222]), .\ootx_payload_o[1][223] (n4568[223]), 
            .\ootx_payload_o[1][224] (n4568[224]), .\ootx_payload_o[1][225] (n4568[225]), 
            .\ootx_payload_o[1][226] (n4568[226]), .\ootx_payload_o[1][227] (n4568[227]), 
            .\ootx_payload_o[1][228] (n4568[228]), .\ootx_payload_o[1][229] (n4568[229]), 
            .\ootx_payload_o[1][230] (n4568[230]), .\ootx_payload_o[1][231] (n4568[231]), 
            .\ootx_payload_o[1][232] (n4568[232]), .\ootx_payload_o[1][233] (n4568[233]), 
            .\ootx_payload_o[1][234] (n4568[234]), .\ootx_payload_o[1][235] (n4568[235]), 
            .\ootx_payload_o[1][236] (n4568[236]), .\ootx_payload_o[1][237] (n4568[237]), 
            .\ootx_payload_o[1][238] (n4568[238]), .\ootx_payload_o[1][239] (n4568[239]), 
            .\ootx_payload_o[1][240] (n4568[240]), .\ootx_payload_o[1][241] (n4568[241]), 
            .\ootx_payload_o[1][242] (n4568[242]), .\ootx_payload_o[1][243] (n4568[243]), 
            .\ootx_payload_o[1][244] (n4568[244]), .\ootx_payload_o[1][245] (n4568[245]), 
            .\ootx_payload_o[1][246] (n4568[246]), .\ootx_payload_o[1][247] (n4568[247]), 
            .\ootx_payload_o[1][248] (n4568[248]), .\ootx_payload_o[1][249] (n4568[249]), 
            .\ootx_payload_o[1][250] (n4568[250]), .\ootx_payload_o[1][251] (n4568[251]), 
            .\ootx_payload_o[1][252] (n4568[252]), .\ootx_payload_o[1][253] (n4568[253]), 
            .\ootx_payload_o[1][254] (n4568[254]), .\ootx_payload_o[1][255] (n4568[255]), 
            .\ootx_payload_o[1][256] (n4568[256]), .\ootx_payload_o[1][257] (n4568[257]), 
            .\ootx_payload_o[1][258] (n4568[258]), .\ootx_payload_o[1][259] (n4568[259]), 
            .\ootx_payload_o[1][260] (n4568[260]), .\ootx_payload_o[1][261] (n4568[261]), 
            .\ootx_payload_o[1][262] (n4568[262]), .\ootx_payload_o[1][263] (n4568[263]), 
            .n860(n860), .n1264(n1264), .ootx_payloads_1_215(ootx_payloads_1_215), 
            .n586(n586), .n1401(n1401), .ootx_payloads_1_214(ootx_payloads_1_214), 
            .n1359(n1359), .ootx_payloads_1_213(ootx_payloads_1_213), .ootx_payloads_1_212(ootx_payloads_1_212), 
            .ootx_payloads_1_211(ootx_payloads_1_211), .n584(n584), .n1402(n1402), 
            .n582(n582), .n1403(n1403), .ootx_payloads_1_210(ootx_payloads_1_210), 
            .n858(n858), .n1265(n1265), .ootx_payloads_1_209(ootx_payloads_1_209), 
            .n580(n580), .n1404(n1404), .ootx_payloads_1_208(ootx_payloads_1_208), 
            .n578(n578), .n1405(n1405), .n972(n972), .n576(n576), .n1406(n1406), 
            .ootx_payloads_1_207(ootx_payloads_1_207), .ootx_payloads_1_206(ootx_payloads_1_206), 
            .ootx_payloads_1_205(ootx_payloads_1_205), .ootx_payloads_1_204(ootx_payloads_1_204), 
            .ootx_payloads_1_203(ootx_payloads_1_203), .n856(n856), .n1266(n1266), 
            .ootx_payloads_1_202(ootx_payloads_1_202), .n574(n574), .n1407(n1407), 
            .n970(n970), .n968(n968), .n572(n572), .n1408(n1408), .ootx_payloads_1_201(ootx_payloads_1_201), 
            .n854(n854), .n1267(n1267), .n570(n570), .n1409(n1409), 
            .n740(n740), .n1324(n1324), .ootx_payloads_1_200(ootx_payloads_1_200), 
            .ootx_payloads_1_199(ootx_payloads_1_199), .n738(n738), .n1325(n1325), 
            .n568(n568), .n1410(n1410), .ootx_payloads_1_198(ootx_payloads_1_198), 
            .n852(n852), .n1268(n1268), .ootx_payloads_1_197(ootx_payloads_1_197), 
            .n566(n566), .n1411(n1411), .ootx_payloads_1_196(ootx_payloads_1_196), 
            .ootx_payloads_1_195(ootx_payloads_1_195), .ootx_payloads_1_194(ootx_payloads_1_194), 
            .ootx_payloads_1_193(ootx_payloads_1_193), .ootx_payloads_1_192(ootx_payloads_1_192), 
            .n564(n564), .n1412(n1412), .n850(n850), .n1269(n1269), 
            .n1360(n1360), .n562(n562), .n1413(n1413), .n708(n708), 
            .n1340(n1340), .n560(n560), .n1414(n1414), .n964(n964), 
            .n9513(n9513), .ootx_payloads_N_1698(ootx_payloads_N_1698), 
            .n558(n558), .n1415(n1415), .ootx_payloads_1_191(ootx_payloads_1_191), 
            .ootx_payloads_1_190(ootx_payloads_1_190), .ootx_payloads_1_189(ootx_payloads_1_189), 
            .ootx_payloads_1_188(ootx_payloads_1_188), .ootx_payloads_1_187(ootx_payloads_1_187), 
            .n848(n848), .n1270(n1270), .ootx_payloads_1_186(ootx_payloads_1_186), 
            .n556(n556), .n1416(n1416), .ootx_payloads_1_185(ootx_payloads_1_185), 
            .ootx_payloads_1_184(ootx_payloads_1_184), .n554(n554), .n1417(n1417), 
            .ootx_payloads_1_183(ootx_payloads_1_183), .n768(n768), .n1310(n1310), 
            .n846(n846), .n1271(n1271), .ootx_payloads_1_182(ootx_payloads_1_182), 
            .n540(n540), .n542(n542), .n544(n544), .n546(n546), .n548(n548), 
            .ootx_payloads_1_181(ootx_payloads_1_181), .n550(n550), .n552(n552), 
            .n1370(n1370), .n736(n736), .n686(n686), .n690(n690), .ootx_payloads_1_180(ootx_payloads_1_180), 
            .n762(n762), .n692(n692), .ootx_payloads_1_179(ootx_payloads_1_179), 
            .n1313(n1313), .n696(n696), .n698(n698), .ootx_payloads_1_178(ootx_payloads_1_178), 
            .n700(n700), .n702(n702), .ootx_payloads_1_177(ootx_payloads_1_177), 
            .n936(n936), .n1226(n1226), .ootx_payloads_1_176(ootx_payloads_1_176), 
            .n704(n704), .ootx_payloads_1_175(ootx_payloads_1_175), .ootx_payloads_1_174(ootx_payloads_1_174), 
            .n706(n706), .ootx_payloads_1_173(ootx_payloads_1_173), .ootx_payloads_1_172(ootx_payloads_1_172), 
            .ootx_payloads_1_171(ootx_payloads_1_171), .ootx_payloads_1_170(ootx_payloads_1_170), 
            .ootx_payloads_1_169(ootx_payloads_1_169), .ootx_payloads_1_168(ootx_payloads_1_168), 
            .ootx_payloads_1_167(ootx_payloads_1_167), .ootx_payloads_1_166(ootx_payloads_1_166), 
            .ootx_payloads_1_165(ootx_payloads_1_165), .n962(n962), .ootx_payloads_1_164(ootx_payloads_1_164), 
            .ootx_payloads_1_163(ootx_payloads_1_163), .ootx_payloads_1_162(ootx_payloads_1_162), 
            .n646(n646), .n1371(n1371), .ootx_payloads_1_161(ootx_payloads_1_161), 
            .ootx_payloads_1_160(ootx_payloads_1_160), .n720(n720), .ootx_payloads_1_159(ootx_payloads_1_159), 
            .n760(n760), .ootx_payloads_1_158(ootx_payloads_1_158), .n1314(n1314), 
            .n642(n642), .n644(n644), .ootx_payloads_1_157(ootx_payloads_1_157), 
            .ootx_payloads_1_156(ootx_payloads_1_156), .ootx_payloads_1_155(ootx_payloads_1_155), 
            .ootx_payloads_1_154(ootx_payloads_1_154), .ootx_payloads_1_153(ootx_payloads_1_153), 
            .ootx_payloads_1_152(ootx_payloads_1_152), .ootx_payloads_1_151(ootx_payloads_1_151), 
            .ootx_payloads_1_150(ootx_payloads_1_150), .ootx_payloads_1_149(ootx_payloads_1_149), 
            .ootx_payloads_1_148(ootx_payloads_1_148), .ootx_payloads_1_147(ootx_payloads_1_147), 
            .n960(n960), .ootx_payloads_1_146(ootx_payloads_1_146), .n770(n770), 
            .n772(n772), .ootx_payloads_1_145(ootx_payloads_1_145), .n774(n774), 
            .n718(n718), .ootx_payloads_1_144(ootx_payloads_1_144), .ootx_payloads_1_143(ootx_payloads_1_143), 
            .n1361(n1361), .n682(n682), .n684(n684), .ootx_payloads_1_142(ootx_payloads_1_142), 
            .n688(n688), .ootx_payloads_1_141(ootx_payloads_1_141), .ootx_payloads_1_140(ootx_payloads_1_140), 
            .n694(n694), .ootx_payloads_1_139(ootx_payloads_1_139), .ootx_payloads_1_138(ootx_payloads_1_138), 
            .ootx_payloads_1_137(ootx_payloads_1_137), .ootx_payloads_1_136(ootx_payloads_1_136), 
            .ootx_payloads_1_135(ootx_payloads_1_135), .n734(n734), .n776(n776), 
            .ootx_payloads_1_134(ootx_payloads_1_134), .ootx_payloads_1_133(ootx_payloads_1_133), 
            .ootx_payloads_1_132(ootx_payloads_1_132), .ootx_payloads_1_131(ootx_payloads_1_131), 
            .n538(n538), .n756(n756), .n758(n758), .ootx_payloads_1_130(ootx_payloads_1_130), 
            .ootx_payloads_1_129(ootx_payloads_1_129), .n728(n728), .ootx_payloads_1_128(ootx_payloads_1_128), 
            .ootx_payloads_1_127(ootx_payloads_1_127), .n714(n714), .n730(n730), 
            .n732(n732), .ootx_payloads_1_126(ootx_payloads_1_126), .ootx_payloads_1_125(ootx_payloads_1_125), 
            .ootx_payloads_1_124(ootx_payloads_1_124), .ootx_payloads_1_123(ootx_payloads_1_123), 
            .ootx_payloads_1_122(ootx_payloads_1_122), .n716(n716), .ootx_payloads_1_121(ootx_payloads_1_121), 
            .ootx_payloads_1_120(ootx_payloads_1_120), .ootx_payloads_1_119(ootx_payloads_1_119), 
            .ootx_payloads_1_118(ootx_payloads_1_118), .ootx_payloads_1_117(ootx_payloads_1_117), 
            .ootx_payloads_1_116(ootx_payloads_1_116), .ootx_payloads_1_115(ootx_payloads_1_115), 
            .n1315(n1315), .ootx_payloads_1_114(ootx_payloads_1_114), .n722(n722), 
            .ootx_payloads_1_113(ootx_payloads_1_113), .ootx_payloads_1_112(ootx_payloads_1_112), 
            .ootx_payloads_1_111(ootx_payloads_1_111), .n1333(n1333), .ootx_payloads_1_110(ootx_payloads_1_110), 
            .n726(n726), .ootx_payloads_1_109(ootx_payloads_1_109), .ootx_payloads_1_108(ootx_payloads_1_108), 
            .ootx_payloads_1_107(ootx_payloads_1_107), .n1418(n1418), .ootx_payloads_1_106(ootx_payloads_1_106), 
            .ootx_payloads_1_105(ootx_payloads_1_105), .ootx_payloads_1_104(ootx_payloads_1_104), 
            .ootx_payloads_1_103(ootx_payloads_1_103), .ootx_payloads_1_102(ootx_payloads_1_102), 
            .ootx_payloads_1_101(ootx_payloads_1_101), .n1216(n1216), .n844(n844), 
            .n1272(n1272), .n1217(n1217), .ootx_payloads_1_100(ootx_payloads_1_100), 
            .n1218(n1218), .ootx_payloads_1_99(ootx_payloads_1_99), .n1219(n1219), 
            .n842(n842), .n1273(n1273), .n1419(n1419), .n1220(n1220), 
            .ootx_payloads_1_98(ootx_payloads_1_98), .ootx_payloads_1_97(ootx_payloads_1_97), 
            .ootx_payloads_1_96(ootx_payloads_1_96), .n1221(n1221), .ootx_payloads_1_95(ootx_payloads_1_95), 
            .ootx_payloads_1_94(ootx_payloads_1_94), .ootx_payloads_1_93(ootx_payloads_1_93), 
            .n1222(n1222), .ootx_payloads_1_92(ootx_payloads_1_92), .n1341(n1341), 
            .ootx_payloads_1_91(ootx_payloads_1_91), .n1223(n1223), .ootx_payloads_1_90(ootx_payloads_1_90), 
            .n1224(n1224), .ootx_payloads_1_89(ootx_payloads_1_89), .ootx_payloads_1_88(ootx_payloads_1_88), 
            .ootx_payloads_1_87(ootx_payloads_1_87), .ootx_payloads_1_86(ootx_payloads_1_86), 
            .n840(n840), .n1274(n1274), .ootx_payloads_1_85(ootx_payloads_1_85), 
            .ootx_payloads_1_84(ootx_payloads_1_84), .ootx_payloads_1_83(ootx_payloads_1_83), 
            .n1420(n1420), .n1227(n1227), .ootx_payloads_1_82(ootx_payloads_1_82), 
            .n1228(n1228), .n838(n838), .n1275(n1275), .ootx_payloads_1_81(ootx_payloads_1_81), 
            .n934(n934), .n1229(n1229), .ootx_payloads_1_80(ootx_payloads_1_80), 
            .ootx_payloads_1_79(ootx_payloads_1_79), .ootx_payloads_1_78(ootx_payloads_1_78), 
            .ootx_payloads_1_77(ootx_payloads_1_77), .ootx_payloads_1_76(ootx_payloads_1_76), 
            .ootx_payloads_1_75(ootx_payloads_1_75), .n1342(n1342), .n1421(n1421), 
            .ootx_payloads_1_74(ootx_payloads_1_74), .n836(n836), .n1276(n1276), 
            .ootx_payloads_1_73(ootx_payloads_1_73), .ootx_payloads_1_72(ootx_payloads_1_72), 
            .n1422(n1422), .n1423(n1423), .n834(n834), .n1277(n1277), 
            .ootx_payloads_1_71(ootx_payloads_1_71), .ootx_payloads_1_70(ootx_payloads_1_70), 
            .n1424(n1424), .ootx_payloads_1_69(ootx_payloads_1_69), .ootx_payloads_1_68(ootx_payloads_1_68), 
            .ootx_payloads_1_67(ootx_payloads_1_67), .ootx_payloads_1_66(ootx_payloads_1_66), 
            .ootx_payloads_1_65(ootx_payloads_1_65), .ootx_payloads_1_64(ootx_payloads_1_64), 
            .n1343(n1343), .n1425(n1425), .ootx_payloads_1_63(ootx_payloads_1_63), 
            .n832(n832), .n1278(n1278), .ootx_payloads_1_62(ootx_payloads_1_62), 
            .ootx_payloads_1_61(ootx_payloads_1_61), .n536(n536), .n1426(n1426), 
            .n1316(n1316), .ootx_payloads_1_60(ootx_payloads_1_60), .n1334(n1334), 
            .ootx_payloads_1_59(ootx_payloads_1_59), .ootx_payloads_1_58(ootx_payloads_1_58), 
            .ootx_payloads_1_57(ootx_payloads_1_57), .n534(n534), .n1427(n1427), 
            .ootx_payloads_1_56(ootx_payloads_1_56), .n830(n830), .n1279(n1279), 
            .n1362(n1362), .ootx_payloads_1_55(ootx_payloads_1_55), .ootx_payloads_1_54(ootx_payloads_1_54), 
            .ootx_payloads_1_53(ootx_payloads_1_53), .n1344(n1344), .n532(n532), 
            .n1428(n1428), .ootx_payloads_1_52(ootx_payloads_1_52), .n828(n828), 
            .n1280(n1280), .n530(n530), .n1429(n1429), .n956(n956), 
            .n1345(n1345), .ootx_payloads_1_51(ootx_payloads_1_51), .ootx_payloads_1_50(ootx_payloads_1_50), 
            .ootx_payloads_1_49(ootx_payloads_1_49), .n954(n954), .n826(n826), 
            .n1281(n1281), .ootx_payloads_1_48(ootx_payloads_1_48), .n528(n528), 
            .n1430(n1430), .ootx_payloads_1_47(ootx_payloads_1_47), .n526(n526), 
            .n1431(n1431), .ootx_payloads_1_46(ootx_payloads_1_46), .ootx_payloads_1_45(ootx_payloads_1_45), 
            .n1346(n1346), .n824(n824), .n1282(n1282), .ootx_payloads_1_44(ootx_payloads_1_44), 
            .n952(n952), .ootx_payloads_1_43(ootx_payloads_1_43), .n524(n524), 
            .n1432(n1432), .\ootx_payloads_N_1730[12] (ootx_payloads_N_1730[12]), 
            .ootx_payloads_1_42(ootx_payloads_1_42), .ootx_payloads_1_41(ootx_payloads_1_41), 
            .ootx_payloads_1_40(ootx_payloads_1_40), .ootx_payloads_1_39(ootx_payloads_1_39), 
            .ootx_payloads_1_38(ootx_payloads_1_38), .ootx_payloads_1_37(ootx_payloads_1_37), 
            .n522(n522), .n1433(n1433), .n822(n822), .n1283(n1283), 
            .n1347(n1347), .n950(n950), .\ootx_payloads_N_1730[11] (ootx_payloads_N_1730[11]), 
            .ootx_payloads_1_36(ootx_payloads_1_36), .ootx_payloads_1_35(ootx_payloads_1_35), 
            .n1326(n1326), .ootx_payloads_1_34(ootx_payloads_1_34), .ootx_payloads_1_33(ootx_payloads_1_33), 
            .n1348(n1348), .n6334(n6334), .ootx_payloads_1_32(ootx_payloads_1_32), 
            .ootx_payloads_1_31(ootx_payloads_1_31), .n51(n51), .n52(n52), 
            .ootx_payloads_1_30(ootx_payloads_1_30), .n948(n948), .\ootx_payloads_N_1730[10] (ootx_payloads_N_1730[10]), 
            .ootx_payloads_1_29(ootx_payloads_1_29), .ootx_payloads_1_28(ootx_payloads_1_28), 
            .n2679(n2679), .n2680(n2680), .n6335(n6335), .n1349(n1349), 
            .ootx_payloads_1_27(ootx_payloads_1_27), .n1317(n1317), .n932(n932), 
            .ootx_payloads_1_26(ootx_payloads_1_26), .n6336(n6336), .n946(n946), 
            .ootx_payloads_1_25(ootx_payloads_1_25), .ootx_payloads_1_24(ootx_payloads_1_24), 
            .ootx_payloads_1_23(ootx_payloads_1_23), .\ootx_payloads_N_1730[9] (ootx_payloads_N_1730[9]), 
            .n1363(n1363), .ootx_payloads_1_22(ootx_payloads_1_22), .n49(n49), 
            .n50(n50), .n9771(n9771), .n820(n820), .n1284(n1284), .ootx_payloads_1_21(ootx_payloads_1_21), 
            .n6337(n6337), .ootx_payloads_1_20(ootx_payloads_1_20), .n1350(n1350), 
            .ootx_payloads_1_19(ootx_payloads_1_19), .ootx_payloads_1_18(ootx_payloads_1_18), 
            .ootx_payloads_1_17(ootx_payloads_1_17), .n944(n944), .n6338(n6338), 
            .ootx_payloads_1_16(ootx_payloads_1_16), .n1351(n1351), .\ootx_payloads_N_1730[8] (ootx_payloads_N_1730[8]), 
            .n47(n47), .n48(n48), .n818(n818), .n1285(n1285), .ootx_payloads_1_15(ootx_payloads_1_15), 
            .ootx_payloads_1_14(ootx_payloads_1_14), .ootx_payloads_1_13(ootx_payloads_1_13), 
            .ootx_payloads_1_12(ootx_payloads_1_12), .n942(n942), .n6339(n6339), 
            .ootx_payloads_1_11(ootx_payloads_1_11), .n45(n45_adj_2271), 
            .n46(n46), .ootx_payloads_1_10(ootx_payloads_1_10), .\ootx_payloads_N_1730[7] (ootx_payloads_N_1730[7]), 
            .n816(n816), .n1286(n1286), .ootx_payloads_1_9(ootx_payloads_1_9), 
            .n6340(n6340), .ootx_payloads_1_8(ootx_payloads_1_8), .crc32s_1_25(crc32s_1_25), 
            .crc32s_1_30(crc32s_1_30), .crc32s_1_27(crc32s_1_27), .crc32s_1_26(crc32s_1_26), 
            .crc32s_1_31(crc32s_1_31), .crc32s_1_29(crc32s_1_29), .crc32s_1_28(crc32s_1_28), 
            .crc32s_1_24(crc32s_1_24), .crc32s_1_23(crc32s_1_23), .crc32s_1_22(crc32s_1_22), 
            .crc32s_1_21(crc32s_1_21), .ootx_payloads_1_7(ootx_payloads_1_7), 
            .crc32s_1_20(crc32s_1_20), .\ootx_payloads_N_1730[6] (ootx_payloads_N_1730[6]), 
            .n1364(n1364), .ootx_payloads_1_6(ootx_payloads_1_6), .ootx_payloads_1_5(ootx_payloads_1_5), 
            .crc32s_1_19(crc32s_1_19), .crc32s_1_18(crc32s_1_18), .crc32s_1_17(crc32s_1_17), 
            .crc32s_1_16(crc32s_1_16), .crc32s_1_15(crc32s_1_15), .n6341(n6341), 
            .crc32s_1_14(crc32s_1_14), .crc32s_1_13(crc32s_1_13), .crc32s_1_12(crc32s_1_12), 
            .crc32s_1_11(crc32s_1_11), .crc32s_1_10(crc32s_1_10), .crc32s_1_9(crc32s_1_9), 
            .crc32s_1_8(crc32s_1_8), .crc32s_1_7(crc32s_1_7), .crc32s_1_6(crc32s_1_6), 
            .crc32s_1_5(crc32s_1_5), .crc32s_1_4(crc32s_1_4), .crc32s_1_3(crc32s_1_3), 
            .crc32s_1_2(crc32s_1_2), .ootx_payloads_1_4(ootx_payloads_1_4), 
            .ootx_payloads_1_3(ootx_payloads_1_3), .crc32s_1_0(crc32s_1_0), 
            .ootx_payloads_1_2(ootx_payloads_1_2), .crc32s_1_1(crc32s_1_1), 
            .\ootx_payloads_N_1730[5] (ootx_payloads_N_1730[5]), .ootx_payloads_1_1(ootx_payloads_1_1), 
            .n43(n43), .n6342(n6342), .n44(n44), .n28(n28_adj_2276), 
            .n814(n814), .n1287(n1287), .n41(n41), .n42(n42), .n1288(n1288), 
            .n1289(n1289), .n1290(n1290), .n1291(n1291), .n1292(n1292), 
            .n1293(n1293), .n1294(n1294), .n1295(n1295), .n1296(n1296), 
            .n1297(n1297), .n1298(n1298), .n1299(n1299), .n1300(n1300), 
            .n1301(n1301), .n1302(n1302), .n1303(n1303), .n1304(n1304), 
            .n1305(n1305), .n1306(n1306), .n1307(n1307), .n1308(n1308), 
            .n1309(n1309), .n1327(n1327), .n1328(n1328), .n1329(n1329), 
            .n1330(n1330), .n1331(n1331), .n1335(n1335), .n1336(n1336), 
            .n1337(n1337), .n1352(n1352), .n1353(n1353), .n1365(n1365), 
            .n1366(n1366), .n1367(n1367), .n1368(n1368), .n1369(n1369), 
            .n1372(n1372), .n1373(n1373), .n11612(n11612), .n3112({n3080, 
            n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
            n3089, n3090, n3091, n3092, n3093_adj_2243, n3094_adj_2244, 
            n3095_adj_2245, n3096_adj_2246, n3097_adj_2247, n3098_adj_2248, 
            n3099_adj_2249, n3100_adj_2250, n3101, n3102, n3103, n3104, 
            n3105, n3106, n3107, n3108, n3109, n3110, n3111}), 
            .n11611(n11611), .n11610(n11610), .n11609(n11609), .n11608(n11608), 
            .n11607(n11607), .n11606(n11606), .n11605(n11605), .n11604(n11604), 
            .n22997(n22997), .n11602(n11602), .n23001(n23001), .n11600(n11600), 
            .n11599(n11599), .n11598(n11598), .n11597(n11597), .n11596(n11596), 
            .n11595(n11595), .n11594(n11594), .n11593(n11593), .n11592(n11592), 
            .n11591(n11591), .n11590(n11590), .n11589(n11589), .n11588(n11588), 
            .n11587(n11587), .n11586(n11586), .n11585(n11585), .n11584(n11584), 
            .n11583(n11583), .n11582(n11582), .n11581(n11581), .n11580(n11580), 
            .n11579(n11579), .n11578(n11578), .n11577(n11577), .n11576(n11576), 
            .n11575(n11575), .n11574(n11574), .n11573(n11573), .n11572(n11572), 
            .n11571(n11571), .n11570(n11570), .n11569(n11569), .n11568(n11568), 
            .n11567(n11567), .n11566(n11566), .n11565(n11565), .n11564(n11564), 
            .n11563(n11563), .n11562(n11562), .n11561(n11561), .n11560(n11560), 
            .n11559(n11559), .n11558(n11558), .n11557(n11557), .n11556(n11556), 
            .n11555(n11555), .n11554(n11554), .n11553(n11553), .n11552(n11552), 
            .n11551(n11551), .n11550(n11550), .n11549(n11549), .n11548(n11548), 
            .n11547(n11547), .n11546(n11546), .n11545(n11545), .n11544(n11544), 
            .n11543(n11543), .n11542(n11542), .n11541(n11541), .n11540(n11540), 
            .n11539(n11539), .n11538(n11538), .n11537(n11537), .n11536(n11536), 
            .n11535(n11535), .n11534(n11534), .n11533(n11533), .n11532(n11532), 
            .n11531(n11531), .n11530(n11530), .n11529(n11529), .n11528(n11528), 
            .n11527(n11527), .n11526(n11526), .n11525(n11525), .n11524(n11524), 
            .n11523(n11523), .n11522(n11522), .n11521(n11521), .n11520(n11520), 
            .n11519(n11519), .n11518(n11518), .n11517(n11517), .n11516(n11516), 
            .n11515(n11515), .n11514(n11514), .n11513(n11513), .n11512(n11512), 
            .n11511(n11511), .n11510(n11510), .n11509(n11509), .n11508(n11508), 
            .n11507(n11507), .n11506(n11506), .n11505(n11505), .n11504(n11504), 
            .n39(n39), .n40(n40), .n812(n812), .n37(n37_adj_2270), .n38(n38), 
            .n6343(n6343), .n810(n810), .n808(n808), .n17(n17), .n19468(n19468), 
            .n806(n806), .n535(n535), .n792(n792), .n804(n804), .n533(n533), 
            .led_c_0(led_c_0), .n790(n790), .led_c_1(led_c_1), .led_c_2(led_c_2), 
            .led_c_3(led_c_3), .led_c_4(led_c_4), .led_c_5(led_c_5), .led_c_6(led_c_6), 
            .n802(n802), .n800(n800), .n531(n531), .n11503(n11503), 
            .n11502(n11502), .n11501(n11501), .n11500(n11500), .n11499(n11499), 
            .n11498(n11498), .n11497(n11497), .n11496(n11496), .n11495(n11495), 
            .n11494(n11494), .n11493(n11493), .n11492(n11492), .n11491(n11491), 
            .n11490(n11490), .n11489(n11489), .n11488(n11488), .n11487(n11487), 
            .n11486(n11486), .n11485(n11485), .n11484(n11484), .n11483(n11483), 
            .n11482(n11482), .n11481(n11481), .n11480(n11480), .n11479(n11479), 
            .n11478(n11478), .n11477(n11477), .n11476(n11476), .n11475(n11475), 
            .n11474(n11474), .n11473(n11473), .n11472(n11472), .n788(n788), 
            .n11471(n11471), .n11470(n11470), .n11469(n11469), .n11468(n11468), 
            .n11467(n11467), .n11466(n11466), .n11465(n11465), .n11464(n11464), 
            .n11463(n11463), .n11462(n11462), .n11461(n11461), .n11460(n11460), 
            .n11459(n11459), .n11458(n11458), .n11457(n11457), .n11456(n11456), 
            .n11455(n11455), .n11454(n11454), .n11453(n11453), .n11452(n11452), 
            .n11451(n11451), .n11450(n11450), .n11449(n11449), .n11448(n11448), 
            .n11447(n11447), .n11446(n11446), .n11445(n11445), .n11444(n11444), 
            .n11443(n11443), .n11442(n11442), .n11441(n11441), .n11440(n11440), 
            .n11439(n11439), .n11438(n11438), .n11437(n11437), .n11436(n11436), 
            .n11435(n11435), .n11434(n11434), .n11433(n11433), .n11432(n11432), 
            .n11431(n11431), .n11430(n11430), .n11429(n11429), .n11428(n11428), 
            .n11427(n11427), .n11426(n11426), .n11425(n11425), .n11424(n11424), 
            .n11423(n11423), .n11422(n11422), .n11421(n11421), .n11420(n11420), 
            .n11419(n11419), .n11418(n11418), .n11417(n11417), .n11416(n11416), 
            .n11415(n11415), .n11414(n11414), .n11413(n11413), .n11412(n11412), 
            .n11411(n11411), .n11410(n11410), .n11409(n11409), .n11408(n11408), 
            .n11407(n11407), .n11406(n11406), .n11405(n11405), .n11404(n11404), 
            .n11403(n11403), .n11402(n11402), .n11401(n11401), .n11400(n11400), 
            .n11399(n11399), .n11398(n11398), .n11397(n11397), .n11396(n11396), 
            .n11395(n11395), .n11394(n11394), .n11393(n11393), .n11392(n11392), 
            .n11391(n11391), .n11390(n11390), .n11389(n11389), .n11388(n11388), 
            .n11387(n11387), .n11386(n11386), .n11385(n11385), .n11384(n11384), 
            .n11383(n11383), .n11382(n11382), .n11381(n11381), .n11380(n11380), 
            .n11379(n11379), .n11378(n11378), .n11377(n11377), .n11376(n11376), 
            .n11375(n11375), .n11374(n11374), .n11373(n11373), .n11372(n11372), 
            .n11371(n11371), .n11370(n11370), .n11369(n11369), .n11368(n11368), 
            .n11367(n11367), .n11366(n11366), .n11365(n11365), .n11364(n11364), 
            .n11363(n11363), .n11362(n11362), .n11361(n11361), .n11360(n11360), 
            .n11359(n11359), .n11358(n11358), .n11357(n11357), .n11356(n11356), 
            .n11355(n11355), .n11354(n11354), .n11353(n11353), .n11352(n11352), 
            .n11351(n11351), .n11350(n11350), .n11349(n11349), .n11348(n11348), 
            .n11347(n11347), .n11346(n11346), .n11345(n11345), .n11344(n11344), 
            .n11343(n11343), .n11342(n11342), .n11341(n11341), .n11340(n11340), 
            .n11339(n11339), .n11338(n11338), .n11337(n11337), .n11336(n11336), 
            .n11335(n11335), .n11334(n11334), .n11333(n11333), .n11332(n11332), 
            .n11331(n11331), .n11330(n11330), .n11329(n11329), .n11328(n11328), 
            .n11327(n11327), .n11326(n11326), .n11325(n11325), .n11324(n11324), 
            .n11323(n11323), .n11322(n11322), .n11321(n11321), .n11320(n11320), 
            .n11319(n11319), .n11318(n11318), .n11317(n11317), .n11316(n11316), 
            .n11315(n11315), .n11314(n11314), .n11313(n11313), .n11312(n11312), 
            .n11311(n11311), .n11310(n11310), .n11309(n11309), .n11308(n11308), 
            .n11307(n11307), .n11306(n11306), .n11305(n11305), .n11304(n11304), 
            .n11303(n11303), .n11302(n11302), .n11301(n11301), .n11300(n11300), 
            .n11299(n11299), .n11298(n11298), .n11297(n11297), .n11296(n11296), 
            .n11295(n11295), .n11294(n11294), .n11293(n11293), .n11292(n11292), 
            .n11291(n11291), .n11290(n11290), .n11289(n11289), .n11288(n11288), 
            .n11287(n11287), .n11286(n11286), .n11285(n11285), .ootx_payloads_1_0(ootx_payloads_1_0), 
            .n6344(n6344), .n798(n798), .n529(n529), .n796(n796), .n6345(n6345), 
            .n786(n786), .n794(n794), .n527(n527), .n6346(n6346), .n784(n784), 
            .n525(n525), .n782(n782), .n523(n523), .n780(n780), .n778(n778), 
            .n521(n521), .n1032(n1032), .\ootx_payloads_N_1730[0] (ootx_payloads_N_1730[0]), 
            .n930(n930), .n940(n940), .sync({sync}), .n1022(n1022), 
            .n1012(n1012), .n1014(n1014), .n1002(n1002), .n1016(n1016), 
            .n1018(n1018), .n1020(n1020), .n1024(n1024), .n1026(n1026), 
            .n1028(n1028), .n1030(n1030), .n11016(n11016), .\ootx_payload_o[0][0] (n4551[0]), 
            .n67(n67), .n65(n65), .n63(n63), .\ootx_states[1][0] (\ootx_states[1] [0]), 
            .n25(n25_adj_2299), .n61(n61), .n59(n59), .n57(n57), .n55(n55), 
            .n53(n53), .n68(n68), .n66(n66), .n64(n64), .n62(n62), 
            .n60(n60), .n58(n58), .n56(n56), .n54(n54_adj_2272), .n20_adj_33(n20_adj_2252), 
            .led_c_7(led_c_7));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(122[25] 134[2])
    SB_LUT4 mux_561_i13_3_lut (.I0(n4568[92]), .I1(n4568[108]), .I2(address_c_0), 
            .I3(GND_net), .O(n4221));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_563_i13_3_lut (.I0(n4568[60]), .I1(n4568[76]), .I2(address_c_0), 
            .I3(GND_net), .O(n4240));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20294_2_lut (.I0(\ootx_crc32_o[0] [11]), .I1(address_c_0), 
            .I2(GND_net), .I3(GND_net), .O(n24662));
    defparam i20294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_475_i12_3_lut (.I0(n4568[11]), .I1(n4568[27]), .I2(address_c_0), 
            .I3(GND_net), .O(n3097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_561_i12_3_lut (.I0(n4568[91]), .I1(n4568[107]), .I2(address_c_0), 
            .I3(GND_net), .O(n4222));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_563_i12_3_lut (.I0(n4568[59]), .I1(n4568[75]), .I2(address_c_0), 
            .I3(GND_net), .O(n4241));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20293_2_lut (.I0(\ootx_crc32_o[0] [10]), .I1(address_c_0), 
            .I2(GND_net), .I3(GND_net), .O(n24661));
    defparam i20293_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_475_i11_3_lut (.I0(n4568[10]), .I1(n4568[26]), .I2(address_c_0), 
            .I3(GND_net), .O(n3098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_561_i11_3_lut (.I0(n4568[90]), .I1(n4568[106]), .I2(address_c_0), 
            .I3(GND_net), .O(n4223));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_563_i11_3_lut (.I0(n4568[58]), .I1(n4568[74]), .I2(address_c_0), 
            .I3(GND_net), .O(n4242));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20306_2_lut (.I0(\ootx_crc32_o[0] [9]), .I1(address_c_0), .I2(GND_net), 
            .I3(GND_net), .O(n24660));
    defparam i20306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_475_i10_3_lut (.I0(n4568[9]), .I1(n4568[25]), .I2(address_c_0), 
            .I3(GND_net), .O(n3099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_561_i10_3_lut (.I0(n4568[89]), .I1(n4568[105]), .I2(address_c_0), 
            .I3(GND_net), .O(n4224));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_563_i10_3_lut (.I0(n4568[57]), .I1(n4568[73]), .I2(address_c_0), 
            .I3(GND_net), .O(n4243));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20274_2_lut (.I0(\ootx_crc32_o[0] [8]), .I1(address_c_0), .I2(GND_net), 
            .I3(GND_net), .O(n24659));
    defparam i20274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_475_i9_3_lut (.I0(n4568[8]), .I1(n4568[24]), .I2(address_c_0), 
            .I3(GND_net), .O(n3100));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_561_i9_3_lut (.I0(n4568[88]), .I1(n4568[104]), .I2(address_c_0), 
            .I3(GND_net), .O(n4225));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_563_i9_3_lut (.I0(n4568[56]), .I1(n4568[72]), .I2(address_c_0), 
            .I3(GND_net), .O(n4244));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20273_4_lut (.I0(\ootx_crc32_o[0] [22]), .I1(n7584), .I2(n4568[38]), 
            .I3(address_c_1), .O(n24658));
    defparam i20273_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12_4_lut (.I0(data_counters_1_15), .I1(n353), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i22_4_lut (.I0(counter_from_last_rise[0]), .I1(n6365), .I2(reset_c), 
            .I3(n2), .O(n8_adj_2280));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i20386_4_lut (.I0(\ootx_crc32_o[0] [19]), .I1(n7584), .I2(n4568[35]), 
            .I3(address_c_1), .O(n24830));
    defparam i20386_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12_4_lut_adj_876 (.I0(data_counters_1_8), .I1(n360), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_876.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_877 (.I0(data_counters_1_14), .I1(n354), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_877.LUT_INIT = 16'haca0;
    SB_DFFER sensor_select__0__i1 (.Q(sensor_select[0]), .C(clock_c), .E(n2208), 
            .D(writedata_c_0), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(103[11] 109[5])
    SB_IO readdata_pad_31 (.PACKAGE_PIN(readdata[31]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_31));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_31.PIN_TYPE = 6'b011001;
    defparam readdata_pad_31.PULLUP = 1'b0;
    defparam readdata_pad_31.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_31.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i12_4_lut_adj_878 (.I0(data_counters_1_13), .I1(n355), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_878.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_879 (.I0(data_counters_1_12), .I1(n356), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23089));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_879.LUT_INIT = 16'haca0;
    SB_LUT4 i1_2_lut (.I0(address_c_1), .I1(address_c_2), .I2(GND_net), 
            .I3(GND_net), .O(n4671));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(address_c_2), .I1(address_c_1), .I2(address_c_0), 
            .I3(GND_net), .O(n4673));
    defparam i1_3_lut.LUT_INIT = 16'h5151;
    SB_LUT4 i1_2_lut_adj_880 (.I0(address_c_1), .I1(address_c_2), .I2(GND_net), 
            .I3(GND_net), .O(n4700));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam i1_2_lut_adj_880.LUT_INIT = 16'h4444;
    SB_IO sensor_signals_pad_0 (.PACKAGE_PIN(sensor_signals[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_0.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_0.PULLUP = 1'b0;
    defparam sensor_signals_pad_0.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i924_3_lut (.I0(address_c_2), .I1(address_c_1), .I2(address_c_0), 
            .I3(GND_net), .O(n4702));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i924_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i12_4_lut_adj_881 (.I0(data_counters_1_11), .I1(n357), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_881.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_882 (.I0(data_counters_1_10), .I1(n358), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_882.LUT_INIT = 16'haca0;
    SB_LUT4 i20317_4_lut (.I0(\ootx_crc32_o[0] [18]), .I1(n7584), .I2(n4568[34]), 
            .I3(address_c_1), .O(n24832));
    defparam i20317_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_557_i16_3_lut (.I0(n4551[95]), .I1(n4551[111]), .I2(address_c_0), 
            .I3(GND_net), .O(n4150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i16_4_lut (.I0(n25726), .I1(n4150), .I2(address_c_2), 
            .I3(address_c_1), .O(n3723));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_557_i15_3_lut (.I0(n4551[94]), .I1(n4551[110]), .I2(address_c_0), 
            .I3(GND_net), .O(n4151));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i15_4_lut (.I0(n25732), .I1(n4151), .I2(address_c_2), 
            .I3(address_c_1), .O(n3724));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_557_i14_3_lut (.I0(n4551[93]), .I1(n4551[109]), .I2(address_c_0), 
            .I3(GND_net), .O(n4152));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i14_4_lut (.I0(n25738), .I1(n4152), .I2(address_c_2), 
            .I3(address_c_1), .O(n3725));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_556_i9_3_lut (.I0(n4551[208]), .I1(n4551[224]), .I2(address_c_0), 
            .I3(GND_net), .O(n4140));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_567_i9_4_lut (.I0(n4140), .I1(n4551[240]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4303));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_553_i9_3_lut (.I0(n4551[136]), .I1(n4551[152]), .I2(address_c_0), 
            .I3(GND_net), .O(n4097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_557_i13_3_lut (.I0(n4551[92]), .I1(n4551[108]), .I2(address_c_0), 
            .I3(GND_net), .O(n4153));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_883 (.I0(data_counters_1_9), .I1(n359), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_883.LUT_INIT = 16'haca0;
    SB_LUT4 mux_529_i13_4_lut (.I0(n25744), .I1(n4153), .I2(address_c_2), 
            .I3(address_c_1), .O(n3726));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_557_i12_3_lut (.I0(n4551[91]), .I1(n4551[107]), .I2(address_c_0), 
            .I3(GND_net), .O(n4154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i12_4_lut (.I0(n25750), .I1(n4154), .I2(address_c_2), 
            .I3(address_c_1), .O(n3727));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_557_i11_3_lut (.I0(n4551[90]), .I1(n4551[106]), .I2(address_c_0), 
            .I3(GND_net), .O(n4155));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i11_4_lut (.I0(n25756), .I1(n4155), .I2(address_c_2), 
            .I3(address_c_1), .O(n3728));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_3_lut_adj_884 (.I0(n13221), .I1(data), .I2(lighthouse[0]), 
            .I3(GND_net), .O(n23974));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i1_3_lut_adj_884.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_2_lut_adj_885 (.I0(data), .I1(n13), .I2(GND_net), .I3(GND_net), 
            .O(n23971));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h4444;
    SB_LUT4 i7175_4_lut (.I0(ootx_payloads_1_0), .I1(data), .I2(n522), 
            .I3(lighthouse[0]), .O(n11285));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7175_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7176_4_lut (.I0(ootx_payloads_1_1), .I1(data), .I2(n524), 
            .I3(lighthouse[0]), .O(n11286));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7176_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7177_4_lut (.I0(ootx_payloads_1_2), .I1(data), .I2(n526), 
            .I3(lighthouse[0]), .O(n11287));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7177_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7178_4_lut (.I0(ootx_payloads_1_3), .I1(data), .I2(n528), 
            .I3(lighthouse[0]), .O(n11288));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7178_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7179_4_lut (.I0(ootx_payloads_1_4), .I1(data), .I2(n530), 
            .I3(lighthouse[0]), .O(n11289));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7179_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7180_4_lut (.I0(ootx_payloads_1_5), .I1(data), .I2(n532), 
            .I3(lighthouse[0]), .O(n11290));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7180_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7181_4_lut (.I0(ootx_payloads_1_6), .I1(data), .I2(n534), 
            .I3(lighthouse[0]), .O(n11291));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7181_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7182_4_lut (.I0(ootx_payloads_1_7), .I1(data), .I2(n536), 
            .I3(lighthouse[0]), .O(n11292));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7182_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7183_4_lut (.I0(ootx_payloads_1_8), .I1(data), .I2(n538), 
            .I3(lighthouse[0]), .O(n11293));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7183_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7184_4_lut (.I0(ootx_payloads_1_9), .I1(data), .I2(n540), 
            .I3(lighthouse[0]), .O(n11294));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7184_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7185_4_lut (.I0(ootx_payloads_1_10), .I1(data), .I2(n542), 
            .I3(lighthouse[0]), .O(n11295));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7185_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7186_4_lut (.I0(ootx_payloads_1_11), .I1(data), .I2(n544), 
            .I3(lighthouse[0]), .O(n11296));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7186_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7187_4_lut (.I0(ootx_payloads_1_12), .I1(data), .I2(n546), 
            .I3(lighthouse[0]), .O(n11297));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7187_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7188_4_lut (.I0(ootx_payloads_1_13), .I1(data), .I2(n548), 
            .I3(lighthouse[0]), .O(n11298));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7188_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7189_4_lut (.I0(ootx_payloads_1_14), .I1(data), .I2(n550), 
            .I3(lighthouse[0]), .O(n11299));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7189_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7190_4_lut (.I0(ootx_payloads_1_15), .I1(data), .I2(n552), 
            .I3(lighthouse[0]), .O(n11300));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7190_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7191_4_lut (.I0(ootx_payloads_1_16), .I1(data), .I2(n554), 
            .I3(lighthouse[0]), .O(n11301));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7191_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7192_4_lut (.I0(ootx_payloads_1_17), .I1(data), .I2(n556), 
            .I3(lighthouse[0]), .O(n11302));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7192_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7193_4_lut (.I0(ootx_payloads_1_18), .I1(data), .I2(n558), 
            .I3(lighthouse[0]), .O(n11303));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7193_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7194_4_lut (.I0(ootx_payloads_1_19), .I1(data), .I2(n560), 
            .I3(lighthouse[0]), .O(n11304));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7194_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7195_4_lut (.I0(ootx_payloads_1_20), .I1(data), .I2(n562), 
            .I3(lighthouse[0]), .O(n11305));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7195_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7196_4_lut (.I0(ootx_payloads_1_21), .I1(data), .I2(n564), 
            .I3(lighthouse[0]), .O(n11306));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7196_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7197_4_lut (.I0(ootx_payloads_1_22), .I1(data), .I2(n566), 
            .I3(lighthouse[0]), .O(n11307));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7197_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7198_4_lut (.I0(ootx_payloads_1_23), .I1(data), .I2(n568), 
            .I3(lighthouse[0]), .O(n11308));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7198_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7199_4_lut (.I0(ootx_payloads_1_24), .I1(data), .I2(n570), 
            .I3(lighthouse[0]), .O(n11309));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7199_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7200_4_lut (.I0(ootx_payloads_1_25), .I1(data), .I2(n572), 
            .I3(lighthouse[0]), .O(n11310));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7200_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7201_4_lut (.I0(ootx_payloads_1_26), .I1(data), .I2(n574), 
            .I3(lighthouse[0]), .O(n11311));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7201_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7202_4_lut (.I0(ootx_payloads_1_27), .I1(data), .I2(n576), 
            .I3(lighthouse[0]), .O(n11312));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7202_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7203_4_lut (.I0(ootx_payloads_1_28), .I1(data), .I2(n578), 
            .I3(lighthouse[0]), .O(n11313));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7203_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7204_4_lut (.I0(ootx_payloads_1_29), .I1(data), .I2(n580), 
            .I3(lighthouse[0]), .O(n11314));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7204_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7205_4_lut (.I0(ootx_payloads_1_30), .I1(data), .I2(n582), 
            .I3(lighthouse[0]), .O(n11315));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7205_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7206_4_lut (.I0(ootx_payloads_1_31), .I1(data), .I2(n584), 
            .I3(lighthouse[0]), .O(n11316));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7206_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7207_4_lut (.I0(ootx_payloads_1_32), .I1(data), .I2(n586), 
            .I3(lighthouse[0]), .O(n11317));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7207_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7208_4_lut (.I0(ootx_payloads_1_33), .I1(data), .I2(n588), 
            .I3(lighthouse[0]), .O(n11318));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7208_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7209_4_lut (.I0(ootx_payloads_1_34), .I1(data), .I2(n590), 
            .I3(lighthouse[0]), .O(n11319));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7209_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7210_4_lut (.I0(ootx_payloads_1_35), .I1(data), .I2(n592), 
            .I3(lighthouse[0]), .O(n11320));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7210_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7211_4_lut (.I0(ootx_payloads_1_36), .I1(data), .I2(n594), 
            .I3(lighthouse[0]), .O(n11321));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7211_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7212_4_lut (.I0(ootx_payloads_1_37), .I1(data), .I2(n596), 
            .I3(lighthouse[0]), .O(n11322));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7212_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7213_4_lut (.I0(ootx_payloads_1_38), .I1(data), .I2(n598), 
            .I3(lighthouse[0]), .O(n11323));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7213_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7214_4_lut (.I0(ootx_payloads_1_39), .I1(data), .I2(n600), 
            .I3(lighthouse[0]), .O(n11324));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7214_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7215_4_lut (.I0(ootx_payloads_1_40), .I1(data), .I2(n602), 
            .I3(lighthouse[0]), .O(n11325));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7215_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7216_4_lut (.I0(ootx_payloads_1_41), .I1(data), .I2(n604), 
            .I3(lighthouse[0]), .O(n11326));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7216_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7217_4_lut (.I0(ootx_payloads_1_42), .I1(data), .I2(n606), 
            .I3(lighthouse[0]), .O(n11327));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7217_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7218_4_lut (.I0(ootx_payloads_1_43), .I1(data), .I2(n608), 
            .I3(lighthouse[0]), .O(n11328));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7218_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7219_4_lut (.I0(ootx_payloads_1_44), .I1(data), .I2(n610), 
            .I3(lighthouse[0]), .O(n11329));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7219_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7220_4_lut (.I0(ootx_payloads_1_45), .I1(data), .I2(n612), 
            .I3(lighthouse[0]), .O(n11330));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7220_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7221_4_lut (.I0(ootx_payloads_1_46), .I1(data), .I2(n614), 
            .I3(lighthouse[0]), .O(n11331));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7221_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7222_4_lut (.I0(ootx_payloads_1_47), .I1(data), .I2(n616), 
            .I3(lighthouse[0]), .O(n11332));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7222_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7223_4_lut (.I0(ootx_payloads_1_48), .I1(data), .I2(n618), 
            .I3(lighthouse[0]), .O(n11333));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7223_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7224_4_lut (.I0(ootx_payloads_1_49), .I1(data), .I2(n620), 
            .I3(lighthouse[0]), .O(n11334));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7224_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7225_4_lut (.I0(ootx_payloads_1_50), .I1(data), .I2(n622), 
            .I3(lighthouse[0]), .O(n11335));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7225_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7226_4_lut (.I0(ootx_payloads_1_51), .I1(data), .I2(n624), 
            .I3(lighthouse[0]), .O(n11336));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7226_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7227_4_lut (.I0(ootx_payloads_1_52), .I1(data), .I2(n626), 
            .I3(lighthouse[0]), .O(n11337));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7227_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7228_4_lut (.I0(ootx_payloads_1_53), .I1(data), .I2(n628), 
            .I3(lighthouse[0]), .O(n11338));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7228_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7229_4_lut (.I0(ootx_payloads_1_54), .I1(data), .I2(n630), 
            .I3(lighthouse[0]), .O(n11339));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7229_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7230_4_lut (.I0(ootx_payloads_1_55), .I1(data), .I2(n632), 
            .I3(lighthouse[0]), .O(n11340));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7230_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7231_4_lut (.I0(ootx_payloads_1_56), .I1(data), .I2(n634), 
            .I3(lighthouse[0]), .O(n11341));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7231_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7232_4_lut (.I0(ootx_payloads_1_57), .I1(data), .I2(n636), 
            .I3(lighthouse[0]), .O(n11342));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7232_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7233_4_lut (.I0(ootx_payloads_1_58), .I1(data), .I2(n638), 
            .I3(lighthouse[0]), .O(n11343));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7233_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7234_4_lut (.I0(ootx_payloads_1_59), .I1(data), .I2(n640), 
            .I3(lighthouse[0]), .O(n11344));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7234_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7235_4_lut (.I0(ootx_payloads_1_60), .I1(data), .I2(n642), 
            .I3(lighthouse[0]), .O(n11345));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7235_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7236_4_lut (.I0(ootx_payloads_1_61), .I1(data), .I2(n644), 
            .I3(lighthouse[0]), .O(n11346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7236_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7237_4_lut (.I0(ootx_payloads_1_62), .I1(data), .I2(n646), 
            .I3(lighthouse[0]), .O(n11347));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7237_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7238_4_lut (.I0(ootx_payloads_1_63), .I1(data), .I2(n648), 
            .I3(lighthouse[0]), .O(n11348));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7238_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7239_4_lut (.I0(ootx_payloads_1_64), .I1(data), .I2(n650), 
            .I3(lighthouse[0]), .O(n11349));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7239_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7240_4_lut (.I0(ootx_payloads_1_65), .I1(data), .I2(n652), 
            .I3(lighthouse[0]), .O(n11350));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7240_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7241_4_lut (.I0(ootx_payloads_1_66), .I1(data), .I2(n654), 
            .I3(lighthouse[0]), .O(n11351));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7241_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7242_4_lut (.I0(ootx_payloads_1_67), .I1(data), .I2(n656), 
            .I3(lighthouse[0]), .O(n11352));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7242_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7243_4_lut (.I0(ootx_payloads_1_68), .I1(data), .I2(n658), 
            .I3(lighthouse[0]), .O(n11353));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7243_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7244_4_lut (.I0(ootx_payloads_1_69), .I1(data), .I2(n660), 
            .I3(lighthouse[0]), .O(n11354));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7244_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7245_4_lut (.I0(ootx_payloads_1_70), .I1(data), .I2(n662), 
            .I3(lighthouse[0]), .O(n11355));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7245_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7246_4_lut (.I0(ootx_payloads_1_71), .I1(data), .I2(n664), 
            .I3(lighthouse[0]), .O(n11356));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7246_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7247_4_lut (.I0(ootx_payloads_1_72), .I1(data), .I2(n666), 
            .I3(lighthouse[0]), .O(n11357));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7247_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7248_4_lut (.I0(ootx_payloads_1_73), .I1(data), .I2(n668), 
            .I3(lighthouse[0]), .O(n11358));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7248_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7249_4_lut (.I0(ootx_payloads_1_74), .I1(data), .I2(n670), 
            .I3(lighthouse[0]), .O(n11359));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7249_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7250_4_lut (.I0(ootx_payloads_1_75), .I1(data), .I2(n672), 
            .I3(lighthouse[0]), .O(n11360));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7250_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7251_4_lut (.I0(ootx_payloads_1_76), .I1(data), .I2(n674), 
            .I3(lighthouse[0]), .O(n11361));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7251_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7252_4_lut (.I0(ootx_payloads_1_77), .I1(data), .I2(n676), 
            .I3(lighthouse[0]), .O(n11362));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7252_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7253_4_lut (.I0(ootx_payloads_1_78), .I1(data), .I2(n678), 
            .I3(lighthouse[0]), .O(n11363));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7253_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7254_4_lut (.I0(ootx_payloads_1_79), .I1(data), .I2(n680), 
            .I3(lighthouse[0]), .O(n11364));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7254_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7255_4_lut (.I0(ootx_payloads_1_80), .I1(data), .I2(n682), 
            .I3(lighthouse[0]), .O(n11365));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7255_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7256_4_lut (.I0(ootx_payloads_1_81), .I1(data), .I2(n684), 
            .I3(lighthouse[0]), .O(n11366));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7256_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7257_4_lut (.I0(ootx_payloads_1_82), .I1(data), .I2(n686), 
            .I3(lighthouse[0]), .O(n11367));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7257_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7258_4_lut (.I0(ootx_payloads_1_83), .I1(data), .I2(n688), 
            .I3(lighthouse[0]), .O(n11368));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7258_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7259_4_lut (.I0(ootx_payloads_1_84), .I1(data), .I2(n690), 
            .I3(lighthouse[0]), .O(n11369));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7259_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7260_4_lut (.I0(ootx_payloads_1_85), .I1(data), .I2(n692), 
            .I3(lighthouse[0]), .O(n11370));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7260_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7261_4_lut (.I0(ootx_payloads_1_86), .I1(data), .I2(n694), 
            .I3(lighthouse[0]), .O(n11371));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7261_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7262_4_lut (.I0(ootx_payloads_1_87), .I1(data), .I2(n696), 
            .I3(lighthouse[0]), .O(n11372));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7262_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7263_4_lut (.I0(ootx_payloads_1_88), .I1(data), .I2(n698), 
            .I3(lighthouse[0]), .O(n11373));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7263_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7264_4_lut (.I0(ootx_payloads_1_89), .I1(data), .I2(n700), 
            .I3(lighthouse[0]), .O(n11374));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7264_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7265_4_lut (.I0(ootx_payloads_1_90), .I1(data), .I2(n702), 
            .I3(lighthouse[0]), .O(n11375));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7265_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7266_4_lut (.I0(ootx_payloads_1_91), .I1(data), .I2(n704), 
            .I3(lighthouse[0]), .O(n11376));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7266_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7267_4_lut (.I0(ootx_payloads_1_92), .I1(data), .I2(n706), 
            .I3(lighthouse[0]), .O(n11377));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7267_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7268_4_lut (.I0(ootx_payloads_1_93), .I1(data), .I2(n708), 
            .I3(lighthouse[0]), .O(n11378));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7268_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7269_4_lut (.I0(ootx_payloads_1_94), .I1(data), .I2(n710), 
            .I3(lighthouse[0]), .O(n11379));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7269_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7270_4_lut (.I0(ootx_payloads_1_95), .I1(data), .I2(n712), 
            .I3(lighthouse[0]), .O(n11380));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7270_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7271_4_lut (.I0(ootx_payloads_1_96), .I1(data), .I2(n714), 
            .I3(lighthouse[0]), .O(n11381));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7271_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7272_4_lut (.I0(ootx_payloads_1_97), .I1(data), .I2(n716), 
            .I3(lighthouse[0]), .O(n11382));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7272_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7273_4_lut (.I0(ootx_payloads_1_98), .I1(data), .I2(n718), 
            .I3(lighthouse[0]), .O(n11383));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7273_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7274_4_lut (.I0(ootx_payloads_1_99), .I1(data), .I2(n720), 
            .I3(lighthouse[0]), .O(n11384));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7274_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7275_4_lut (.I0(ootx_payloads_1_100), .I1(data), .I2(n722), 
            .I3(lighthouse[0]), .O(n11385));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7275_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7276_4_lut (.I0(ootx_payloads_1_101), .I1(data), .I2(n724), 
            .I3(lighthouse[0]), .O(n11386));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7276_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7277_4_lut (.I0(ootx_payloads_1_102), .I1(data), .I2(n726), 
            .I3(lighthouse[0]), .O(n11387));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7277_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7278_4_lut (.I0(ootx_payloads_1_103), .I1(data), .I2(n728), 
            .I3(lighthouse[0]), .O(n11388));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7278_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7279_4_lut (.I0(ootx_payloads_1_104), .I1(data), .I2(n730), 
            .I3(lighthouse[0]), .O(n11389));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7279_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7280_4_lut (.I0(ootx_payloads_1_105), .I1(data), .I2(n732), 
            .I3(lighthouse[0]), .O(n11390));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7280_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7281_4_lut (.I0(ootx_payloads_1_106), .I1(data), .I2(n734), 
            .I3(lighthouse[0]), .O(n11391));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7281_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7282_4_lut (.I0(ootx_payloads_1_107), .I1(data), .I2(n736), 
            .I3(lighthouse[0]), .O(n11392));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7282_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7283_4_lut (.I0(ootx_payloads_1_108), .I1(data), .I2(n738), 
            .I3(lighthouse[0]), .O(n11393));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7283_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7284_4_lut (.I0(ootx_payloads_1_109), .I1(data), .I2(n740), 
            .I3(lighthouse[0]), .O(n11394));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7284_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7285_4_lut (.I0(ootx_payloads_1_110), .I1(data), .I2(n742), 
            .I3(lighthouse[0]), .O(n11395));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7285_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7286_4_lut (.I0(ootx_payloads_1_111), .I1(data), .I2(n744), 
            .I3(lighthouse[0]), .O(n11396));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7286_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7287_4_lut (.I0(ootx_payloads_1_112), .I1(data), .I2(n746), 
            .I3(lighthouse[0]), .O(n11397));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7287_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7288_4_lut (.I0(ootx_payloads_1_113), .I1(data), .I2(n748), 
            .I3(lighthouse[0]), .O(n11398));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7288_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7289_4_lut (.I0(ootx_payloads_1_114), .I1(data), .I2(n750), 
            .I3(lighthouse[0]), .O(n11399));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7289_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7290_4_lut (.I0(ootx_payloads_1_115), .I1(data), .I2(n752), 
            .I3(lighthouse[0]), .O(n11400));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7290_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7291_4_lut (.I0(ootx_payloads_1_116), .I1(data), .I2(n754), 
            .I3(lighthouse[0]), .O(n11401));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7291_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7292_4_lut (.I0(ootx_payloads_1_117), .I1(data), .I2(n756), 
            .I3(lighthouse[0]), .O(n11402));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7292_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7293_4_lut (.I0(ootx_payloads_1_118), .I1(data), .I2(n758), 
            .I3(lighthouse[0]), .O(n11403));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7293_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7294_4_lut (.I0(ootx_payloads_1_119), .I1(data), .I2(n760), 
            .I3(lighthouse[0]), .O(n11404));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7294_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7295_4_lut (.I0(ootx_payloads_1_120), .I1(data), .I2(n762), 
            .I3(lighthouse[0]), .O(n11405));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7295_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7296_4_lut (.I0(ootx_payloads_1_121), .I1(data), .I2(n764), 
            .I3(lighthouse[0]), .O(n11406));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7296_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7297_4_lut (.I0(ootx_payloads_1_122), .I1(data), .I2(n766), 
            .I3(lighthouse[0]), .O(n11407));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7297_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7298_4_lut (.I0(ootx_payloads_1_123), .I1(data), .I2(n768), 
            .I3(lighthouse[0]), .O(n11408));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7298_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7299_4_lut (.I0(ootx_payloads_1_124), .I1(data), .I2(n770), 
            .I3(lighthouse[0]), .O(n11409));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7299_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7300_4_lut (.I0(ootx_payloads_1_125), .I1(data), .I2(n772), 
            .I3(lighthouse[0]), .O(n11410));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7300_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7301_4_lut (.I0(ootx_payloads_1_126), .I1(data), .I2(n774), 
            .I3(lighthouse[0]), .O(n11411));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7301_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7302_4_lut (.I0(ootx_payloads_1_127), .I1(data), .I2(n776), 
            .I3(lighthouse[0]), .O(n11412));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7302_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7303_4_lut (.I0(ootx_payloads_1_128), .I1(data), .I2(n778), 
            .I3(lighthouse[0]), .O(n11413));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7303_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7304_4_lut (.I0(ootx_payloads_1_129), .I1(data), .I2(n780), 
            .I3(lighthouse[0]), .O(n11414));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7304_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7305_4_lut (.I0(ootx_payloads_1_130), .I1(data), .I2(n782), 
            .I3(lighthouse[0]), .O(n11415));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7305_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7306_4_lut (.I0(ootx_payloads_1_131), .I1(data), .I2(n784), 
            .I3(lighthouse[0]), .O(n11416));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7306_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7307_4_lut (.I0(ootx_payloads_1_132), .I1(data), .I2(n786), 
            .I3(lighthouse[0]), .O(n11417));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7307_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7308_4_lut (.I0(ootx_payloads_1_133), .I1(data), .I2(n788), 
            .I3(lighthouse[0]), .O(n11418));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7308_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7309_4_lut (.I0(ootx_payloads_1_134), .I1(data), .I2(n790), 
            .I3(lighthouse[0]), .O(n11419));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7309_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7310_4_lut (.I0(ootx_payloads_1_135), .I1(data), .I2(n792), 
            .I3(lighthouse[0]), .O(n11420));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7310_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7311_4_lut (.I0(ootx_payloads_1_136), .I1(data), .I2(n794), 
            .I3(lighthouse[0]), .O(n11421));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7311_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7312_4_lut (.I0(ootx_payloads_1_137), .I1(data), .I2(n796), 
            .I3(lighthouse[0]), .O(n11422));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7312_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7313_4_lut (.I0(ootx_payloads_1_138), .I1(data), .I2(n798), 
            .I3(lighthouse[0]), .O(n11423));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7313_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7314_4_lut (.I0(ootx_payloads_1_139), .I1(data), .I2(n800), 
            .I3(lighthouse[0]), .O(n11424));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7314_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7315_4_lut (.I0(ootx_payloads_1_140), .I1(data), .I2(n802), 
            .I3(lighthouse[0]), .O(n11425));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7315_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7316_4_lut (.I0(ootx_payloads_1_141), .I1(data), .I2(n804), 
            .I3(lighthouse[0]), .O(n11426));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7316_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7317_4_lut (.I0(ootx_payloads_1_142), .I1(data), .I2(n806), 
            .I3(lighthouse[0]), .O(n11427));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7317_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7318_4_lut (.I0(ootx_payloads_1_143), .I1(data), .I2(n808), 
            .I3(lighthouse[0]), .O(n11428));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7318_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7319_4_lut (.I0(ootx_payloads_1_144), .I1(data), .I2(n810), 
            .I3(lighthouse[0]), .O(n11429));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7319_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7320_4_lut (.I0(ootx_payloads_1_145), .I1(data), .I2(n812), 
            .I3(lighthouse[0]), .O(n11430));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7320_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7321_4_lut (.I0(ootx_payloads_1_146), .I1(data), .I2(n814), 
            .I3(lighthouse[0]), .O(n11431));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7321_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7322_4_lut (.I0(ootx_payloads_1_147), .I1(data), .I2(n816), 
            .I3(lighthouse[0]), .O(n11432));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7322_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7323_4_lut (.I0(ootx_payloads_1_148), .I1(data), .I2(n818), 
            .I3(lighthouse[0]), .O(n11433));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7323_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7324_4_lut (.I0(ootx_payloads_1_149), .I1(data), .I2(n820), 
            .I3(lighthouse[0]), .O(n11434));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7324_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7325_4_lut (.I0(ootx_payloads_1_150), .I1(data), .I2(n822), 
            .I3(lighthouse[0]), .O(n11435));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7325_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7326_4_lut (.I0(ootx_payloads_1_151), .I1(data), .I2(n824), 
            .I3(lighthouse[0]), .O(n11436));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7326_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7327_4_lut (.I0(ootx_payloads_1_152), .I1(data), .I2(n826), 
            .I3(lighthouse[0]), .O(n11437));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7327_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7328_4_lut (.I0(ootx_payloads_1_153), .I1(data), .I2(n828), 
            .I3(lighthouse[0]), .O(n11438));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7328_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7329_4_lut (.I0(ootx_payloads_1_154), .I1(data), .I2(n830), 
            .I3(lighthouse[0]), .O(n11439));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7329_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7330_4_lut (.I0(ootx_payloads_1_155), .I1(data), .I2(n832), 
            .I3(lighthouse[0]), .O(n11440));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7330_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7331_4_lut (.I0(ootx_payloads_1_156), .I1(data), .I2(n834), 
            .I3(lighthouse[0]), .O(n11441));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7331_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7332_4_lut (.I0(ootx_payloads_1_157), .I1(data), .I2(n836), 
            .I3(lighthouse[0]), .O(n11442));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7332_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7333_4_lut (.I0(ootx_payloads_1_158), .I1(data), .I2(n838), 
            .I3(lighthouse[0]), .O(n11443));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7333_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7334_4_lut (.I0(ootx_payloads_1_159), .I1(data), .I2(n840), 
            .I3(lighthouse[0]), .O(n11444));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7334_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7335_4_lut (.I0(ootx_payloads_1_160), .I1(data), .I2(n842), 
            .I3(lighthouse[0]), .O(n11445));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7335_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7336_4_lut (.I0(ootx_payloads_1_161), .I1(data), .I2(n844), 
            .I3(lighthouse[0]), .O(n11446));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7336_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7337_4_lut (.I0(ootx_payloads_1_162), .I1(data), .I2(n846), 
            .I3(lighthouse[0]), .O(n11447));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7337_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7338_4_lut (.I0(ootx_payloads_1_163), .I1(data), .I2(n848), 
            .I3(lighthouse[0]), .O(n11448));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7338_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7339_4_lut (.I0(ootx_payloads_1_164), .I1(data), .I2(n850), 
            .I3(lighthouse[0]), .O(n11449));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7339_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7340_4_lut (.I0(ootx_payloads_1_165), .I1(data), .I2(n852), 
            .I3(lighthouse[0]), .O(n11450));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7340_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7341_4_lut (.I0(ootx_payloads_1_166), .I1(data), .I2(n854), 
            .I3(lighthouse[0]), .O(n11451));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7341_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7342_4_lut (.I0(ootx_payloads_1_167), .I1(data), .I2(n856), 
            .I3(lighthouse[0]), .O(n11452));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7342_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7343_4_lut (.I0(ootx_payloads_1_168), .I1(data), .I2(n858), 
            .I3(lighthouse[0]), .O(n11453));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7343_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7344_4_lut (.I0(ootx_payloads_1_169), .I1(data), .I2(n860), 
            .I3(lighthouse[0]), .O(n11454));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7344_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7345_4_lut (.I0(ootx_payloads_1_170), .I1(data), .I2(n862), 
            .I3(lighthouse[0]), .O(n11455));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7345_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7346_4_lut (.I0(ootx_payloads_1_171), .I1(data), .I2(n864), 
            .I3(lighthouse[0]), .O(n11456));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7346_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7347_4_lut (.I0(ootx_payloads_1_172), .I1(data), .I2(n866), 
            .I3(lighthouse[0]), .O(n11457));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7347_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7348_4_lut (.I0(ootx_payloads_1_173), .I1(data), .I2(n868), 
            .I3(lighthouse[0]), .O(n11458));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7348_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7349_4_lut (.I0(ootx_payloads_1_174), .I1(data), .I2(n870), 
            .I3(lighthouse[0]), .O(n11459));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7349_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7350_4_lut (.I0(ootx_payloads_1_175), .I1(data), .I2(n872), 
            .I3(lighthouse[0]), .O(n11460));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7350_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7351_4_lut (.I0(ootx_payloads_1_176), .I1(data), .I2(n874), 
            .I3(lighthouse[0]), .O(n11461));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7351_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7352_4_lut (.I0(ootx_payloads_1_177), .I1(data), .I2(n876), 
            .I3(lighthouse[0]), .O(n11462));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7352_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7353_4_lut (.I0(ootx_payloads_1_178), .I1(data), .I2(n878), 
            .I3(lighthouse[0]), .O(n11463));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7353_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7354_4_lut (.I0(ootx_payloads_1_179), .I1(data), .I2(n880), 
            .I3(lighthouse[0]), .O(n11464));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7354_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7355_4_lut (.I0(ootx_payloads_1_180), .I1(data), .I2(n882), 
            .I3(lighthouse[0]), .O(n11465));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7355_4_lut.LUT_INIT = 16'hcaaa;
    SB_IO readdata_pad_30 (.PACKAGE_PIN(readdata[30]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_30));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_30.PIN_TYPE = 6'b011001;
    defparam readdata_pad_30.PULLUP = 1'b0;
    defparam readdata_pad_30.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_30.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_1 (.PACKAGE_PIN(sensor_signals[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_1));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_1.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_1.PULLUP = 1'b0;
    defparam sensor_signals_pad_1.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_2 (.PACKAGE_PIN(sensor_signals[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_2));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_2.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_2.PULLUP = 1'b0;
    defparam sensor_signals_pad_2.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_3 (.PACKAGE_PIN(sensor_signals[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_3));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_3.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_3.PULLUP = 1'b0;
    defparam sensor_signals_pad_3.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_4 (.PACKAGE_PIN(sensor_signals[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_4));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_4.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_4.PULLUP = 1'b0;
    defparam sensor_signals_pad_4.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_5 (.PACKAGE_PIN(sensor_signals[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_5));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_5.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_5.PULLUP = 1'b0;
    defparam sensor_signals_pad_5.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_6 (.PACKAGE_PIN(sensor_signals[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_6));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_6.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_6.PULLUP = 1'b0;
    defparam sensor_signals_pad_6.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO sensor_signals_pad_7 (.PACKAGE_PIN(sensor_signals[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(sensor_signals_c_7));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sensor_signals_pad_7.PIN_TYPE = 6'b000001;
    defparam sensor_signals_pad_7.PULLUP = 1'b0;
    defparam sensor_signals_pad_7.NEG_TRIGGER = 1'b0;
    defparam sensor_signals_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_0 (.PACKAGE_PIN(writedata[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_0.PIN_TYPE = 6'b000001;
    defparam writedata_pad_0.PULLUP = 1'b0;
    defparam writedata_pad_0.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_1 (.PACKAGE_PIN(writedata[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_1));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_1.PIN_TYPE = 6'b000001;
    defparam writedata_pad_1.PULLUP = 1'b0;
    defparam writedata_pad_1.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_2 (.PACKAGE_PIN(writedata[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_2));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_2.PIN_TYPE = 6'b000001;
    defparam writedata_pad_2.PULLUP = 1'b0;
    defparam writedata_pad_2.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_3 (.PACKAGE_PIN(writedata[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_3));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_3.PIN_TYPE = 6'b000001;
    defparam writedata_pad_3.PULLUP = 1'b0;
    defparam writedata_pad_3.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_4 (.PACKAGE_PIN(writedata[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_4));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_4.PIN_TYPE = 6'b000001;
    defparam writedata_pad_4.PULLUP = 1'b0;
    defparam writedata_pad_4.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_5 (.PACKAGE_PIN(writedata[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_5));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_5.PIN_TYPE = 6'b000001;
    defparam writedata_pad_5.PULLUP = 1'b0;
    defparam writedata_pad_5.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_6 (.PACKAGE_PIN(writedata[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_6));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_6.PIN_TYPE = 6'b000001;
    defparam writedata_pad_6.PULLUP = 1'b0;
    defparam writedata_pad_6.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_7 (.PACKAGE_PIN(writedata[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_7));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_7.PIN_TYPE = 6'b000001;
    defparam writedata_pad_7.PULLUP = 1'b0;
    defparam writedata_pad_7.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_8 (.PACKAGE_PIN(writedata[8]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_8));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_8.PIN_TYPE = 6'b000001;
    defparam writedata_pad_8.PULLUP = 1'b0;
    defparam writedata_pad_8.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_8.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_9 (.PACKAGE_PIN(writedata[9]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_9));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_9.PIN_TYPE = 6'b000001;
    defparam writedata_pad_9.PULLUP = 1'b0;
    defparam writedata_pad_9.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_9.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_10 (.PACKAGE_PIN(writedata[10]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_10));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_10.PIN_TYPE = 6'b000001;
    defparam writedata_pad_10.PULLUP = 1'b0;
    defparam writedata_pad_10.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_10.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_11 (.PACKAGE_PIN(writedata[11]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_11));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_11.PIN_TYPE = 6'b000001;
    defparam writedata_pad_11.PULLUP = 1'b0;
    defparam writedata_pad_11.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_11.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_12 (.PACKAGE_PIN(writedata[12]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_12));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_12.PIN_TYPE = 6'b000001;
    defparam writedata_pad_12.PULLUP = 1'b0;
    defparam writedata_pad_12.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_12.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_13 (.PACKAGE_PIN(writedata[13]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_13));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_13.PIN_TYPE = 6'b000001;
    defparam writedata_pad_13.PULLUP = 1'b0;
    defparam writedata_pad_13.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_13.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_14 (.PACKAGE_PIN(writedata[14]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_14));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_14.PIN_TYPE = 6'b000001;
    defparam writedata_pad_14.PULLUP = 1'b0;
    defparam writedata_pad_14.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_14.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_15 (.PACKAGE_PIN(writedata[15]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_15));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_15.PIN_TYPE = 6'b000001;
    defparam writedata_pad_15.PULLUP = 1'b0;
    defparam writedata_pad_15.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_15.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_16 (.PACKAGE_PIN(writedata[16]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_16));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_16.PIN_TYPE = 6'b000001;
    defparam writedata_pad_16.PULLUP = 1'b0;
    defparam writedata_pad_16.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_16.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_17 (.PACKAGE_PIN(writedata[17]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_17));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_17.PIN_TYPE = 6'b000001;
    defparam writedata_pad_17.PULLUP = 1'b0;
    defparam writedata_pad_17.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_17.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_18 (.PACKAGE_PIN(writedata[18]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_18));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_18.PIN_TYPE = 6'b000001;
    defparam writedata_pad_18.PULLUP = 1'b0;
    defparam writedata_pad_18.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_18.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_19 (.PACKAGE_PIN(writedata[19]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_19));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_19.PIN_TYPE = 6'b000001;
    defparam writedata_pad_19.PULLUP = 1'b0;
    defparam writedata_pad_19.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_19.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_20 (.PACKAGE_PIN(writedata[20]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_20));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_20.PIN_TYPE = 6'b000001;
    defparam writedata_pad_20.PULLUP = 1'b0;
    defparam writedata_pad_20.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_20.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_21 (.PACKAGE_PIN(writedata[21]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_21));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_21.PIN_TYPE = 6'b000001;
    defparam writedata_pad_21.PULLUP = 1'b0;
    defparam writedata_pad_21.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_21.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_22 (.PACKAGE_PIN(writedata[22]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_22));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_22.PIN_TYPE = 6'b000001;
    defparam writedata_pad_22.PULLUP = 1'b0;
    defparam writedata_pad_22.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_22.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_23 (.PACKAGE_PIN(writedata[23]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_23));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_23.PIN_TYPE = 6'b000001;
    defparam writedata_pad_23.PULLUP = 1'b0;
    defparam writedata_pad_23.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_23.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_24 (.PACKAGE_PIN(writedata[24]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_24));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_24.PIN_TYPE = 6'b000001;
    defparam writedata_pad_24.PULLUP = 1'b0;
    defparam writedata_pad_24.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_24.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_25 (.PACKAGE_PIN(writedata[25]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_25));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_25.PIN_TYPE = 6'b000001;
    defparam writedata_pad_25.PULLUP = 1'b0;
    defparam writedata_pad_25.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_25.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_26 (.PACKAGE_PIN(writedata[26]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_26));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_26.PIN_TYPE = 6'b000001;
    defparam writedata_pad_26.PULLUP = 1'b0;
    defparam writedata_pad_26.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_26.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_27 (.PACKAGE_PIN(writedata[27]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_27));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_27.PIN_TYPE = 6'b000001;
    defparam writedata_pad_27.PULLUP = 1'b0;
    defparam writedata_pad_27.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_27.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_28 (.PACKAGE_PIN(writedata[28]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_28));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_28.PIN_TYPE = 6'b000001;
    defparam writedata_pad_28.PULLUP = 1'b0;
    defparam writedata_pad_28.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_28.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_29 (.PACKAGE_PIN(writedata[29]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_29));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_29.PIN_TYPE = 6'b000001;
    defparam writedata_pad_29.PULLUP = 1'b0;
    defparam writedata_pad_29.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_29.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_30 (.PACKAGE_PIN(writedata[30]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_30));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_30.PIN_TYPE = 6'b000001;
    defparam writedata_pad_30.PULLUP = 1'b0;
    defparam writedata_pad_30.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_30.IO_STANDARD = "SB_LVCMOS";
    SB_IO writedata_pad_31 (.PACKAGE_PIN(writedata[31]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(writedata_c_31));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam writedata_pad_31.PIN_TYPE = 6'b000001;
    defparam writedata_pad_31.PULLUP = 1'b0;
    defparam writedata_pad_31.NEG_TRIGGER = 1'b0;
    defparam writedata_pad_31.IO_STANDARD = "SB_LVCMOS";
    SB_IO write_pad (.PACKAGE_PIN(write), .OUTPUT_ENABLE(VCC_net), .D_IN_0(write_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam write_pad.PIN_TYPE = 6'b000001;
    defparam write_pad.PULLUP = 1'b0;
    defparam write_pad.NEG_TRIGGER = 1'b0;
    defparam write_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO address_pad_0 (.PACKAGE_PIN(address[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(address_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam address_pad_0.PIN_TYPE = 6'b000001;
    defparam address_pad_0.PULLUP = 1'b0;
    defparam address_pad_0.NEG_TRIGGER = 1'b0;
    defparam address_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO address_pad_1 (.PACKAGE_PIN(address[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(address_c_1));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam address_pad_1.PIN_TYPE = 6'b000001;
    defparam address_pad_1.PULLUP = 1'b0;
    defparam address_pad_1.NEG_TRIGGER = 1'b0;
    defparam address_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO address_pad_2 (.PACKAGE_PIN(address[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(address_c_2));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam address_pad_2.PIN_TYPE = 6'b000001;
    defparam address_pad_2.PULLUP = 1'b0;
    defparam address_pad_2.NEG_TRIGGER = 1'b0;
    defparam address_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO address_pad_3 (.PACKAGE_PIN(address[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(address_c_3));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam address_pad_3.PIN_TYPE = 6'b000001;
    defparam address_pad_3.PULLUP = 1'b0;
    defparam address_pad_3.NEG_TRIGGER = 1'b0;
    defparam address_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO address_pad_4 (.PACKAGE_PIN(address[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(address_c_4));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam address_pad_4.PIN_TYPE = 6'b000001;
    defparam address_pad_4.PULLUP = 1'b0;
    defparam address_pad_4.NEG_TRIGGER = 1'b0;
    defparam address_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO address_pad_5 (.PACKAGE_PIN(address[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(address_c_5));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam address_pad_5.PIN_TYPE = 6'b000001;
    defparam address_pad_5.PULLUP = 1'b0;
    defparam address_pad_5.NEG_TRIGGER = 1'b0;
    defparam address_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO reset_pad (.PACKAGE_PIN(reset), .OUTPUT_ENABLE(VCC_net), .D_IN_0(reset_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam reset_pad.PIN_TYPE = 6'b000001;
    defparam reset_pad.PULLUP = 1'b0;
    defparam reset_pad.NEG_TRIGGER = 1'b0;
    defparam reset_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO clock_pad (.PACKAGE_PIN(clock), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clock_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(40[8:13])
    defparam clock_pad.PIN_TYPE = 6'b000001;
    defparam clock_pad.PULLUP = 1'b0;
    defparam clock_pad.NEG_TRIGGER = 1'b0;
    defparam clock_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_0 (.PACKAGE_PIN(led[0]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_0.PIN_TYPE = 6'b011001;
    defparam led_pad_0.PULLUP = 1'b0;
    defparam led_pad_0.NEG_TRIGGER = 1'b0;
    defparam led_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_1 (.PACKAGE_PIN(led[1]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_1));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_1.PIN_TYPE = 6'b011001;
    defparam led_pad_1.PULLUP = 1'b0;
    defparam led_pad_1.NEG_TRIGGER = 1'b0;
    defparam led_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_2 (.PACKAGE_PIN(led[2]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_2));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_2.PIN_TYPE = 6'b011001;
    defparam led_pad_2.PULLUP = 1'b0;
    defparam led_pad_2.NEG_TRIGGER = 1'b0;
    defparam led_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_3 (.PACKAGE_PIN(led[3]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_3));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_3.PIN_TYPE = 6'b011001;
    defparam led_pad_3.PULLUP = 1'b0;
    defparam led_pad_3.NEG_TRIGGER = 1'b0;
    defparam led_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_4 (.PACKAGE_PIN(led[4]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_4));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_4.PIN_TYPE = 6'b011001;
    defparam led_pad_4.PULLUP = 1'b0;
    defparam led_pad_4.NEG_TRIGGER = 1'b0;
    defparam led_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_5 (.PACKAGE_PIN(led[5]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_5));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_5.PIN_TYPE = 6'b011001;
    defparam led_pad_5.PULLUP = 1'b0;
    defparam led_pad_5.NEG_TRIGGER = 1'b0;
    defparam led_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_6 (.PACKAGE_PIN(led[6]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_6));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_6.PIN_TYPE = 6'b011001;
    defparam led_pad_6.PULLUP = 1'b0;
    defparam led_pad_6.NEG_TRIGGER = 1'b0;
    defparam led_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO led_pad_7 (.PACKAGE_PIN(led[7]), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(led_c_7));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam led_pad_7.PIN_TYPE = 6'b011001;
    defparam led_pad_7.PULLUP = 1'b0;
    defparam led_pad_7.NEG_TRIGGER = 1'b0;
    defparam led_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO uart_tx_pad (.PACKAGE_PIN(uart_tx), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam uart_tx_pad.PIN_TYPE = 6'b011001;
    defparam uart_tx_pad.PULLUP = 1'b0;
    defparam uart_tx_pad.NEG_TRIGGER = 1'b0;
    defparam uart_tx_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO waitrequest_pad (.PACKAGE_PIN(waitrequest), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(waitrequest_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam waitrequest_pad.PIN_TYPE = 6'b011001;
    defparam waitrequest_pad.PULLUP = 1'b0;
    defparam waitrequest_pad.NEG_TRIGGER = 1'b0;
    defparam waitrequest_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_0 (.PACKAGE_PIN(readdata[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_0.PIN_TYPE = 6'b011001;
    defparam readdata_pad_0.PULLUP = 1'b0;
    defparam readdata_pad_0.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_1 (.PACKAGE_PIN(readdata[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_1));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_1.PIN_TYPE = 6'b011001;
    defparam readdata_pad_1.PULLUP = 1'b0;
    defparam readdata_pad_1.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_2 (.PACKAGE_PIN(readdata[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_2));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_2.PIN_TYPE = 6'b011001;
    defparam readdata_pad_2.PULLUP = 1'b0;
    defparam readdata_pad_2.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_3 (.PACKAGE_PIN(readdata[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_3));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_3.PIN_TYPE = 6'b011001;
    defparam readdata_pad_3.PULLUP = 1'b0;
    defparam readdata_pad_3.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_4 (.PACKAGE_PIN(readdata[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_4));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_4.PIN_TYPE = 6'b011001;
    defparam readdata_pad_4.PULLUP = 1'b0;
    defparam readdata_pad_4.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_5 (.PACKAGE_PIN(readdata[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_5));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_5.PIN_TYPE = 6'b011001;
    defparam readdata_pad_5.PULLUP = 1'b0;
    defparam readdata_pad_5.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_6 (.PACKAGE_PIN(readdata[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_6));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_6.PIN_TYPE = 6'b011001;
    defparam readdata_pad_6.PULLUP = 1'b0;
    defparam readdata_pad_6.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_7 (.PACKAGE_PIN(readdata[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_7));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_7.PIN_TYPE = 6'b011001;
    defparam readdata_pad_7.PULLUP = 1'b0;
    defparam readdata_pad_7.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_8 (.PACKAGE_PIN(readdata[8]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_8));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_8.PIN_TYPE = 6'b011001;
    defparam readdata_pad_8.PULLUP = 1'b0;
    defparam readdata_pad_8.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_8.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_9 (.PACKAGE_PIN(readdata[9]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_9));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_9.PIN_TYPE = 6'b011001;
    defparam readdata_pad_9.PULLUP = 1'b0;
    defparam readdata_pad_9.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_9.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_10 (.PACKAGE_PIN(readdata[10]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_10));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_10.PIN_TYPE = 6'b011001;
    defparam readdata_pad_10.PULLUP = 1'b0;
    defparam readdata_pad_10.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_10.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_11 (.PACKAGE_PIN(readdata[11]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_11));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_11.PIN_TYPE = 6'b011001;
    defparam readdata_pad_11.PULLUP = 1'b0;
    defparam readdata_pad_11.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_11.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_12 (.PACKAGE_PIN(readdata[12]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_12));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_12.PIN_TYPE = 6'b011001;
    defparam readdata_pad_12.PULLUP = 1'b0;
    defparam readdata_pad_12.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_12.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_13 (.PACKAGE_PIN(readdata[13]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_13));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_13.PIN_TYPE = 6'b011001;
    defparam readdata_pad_13.PULLUP = 1'b0;
    defparam readdata_pad_13.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_13.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_14 (.PACKAGE_PIN(readdata[14]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_14));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_14.PIN_TYPE = 6'b011001;
    defparam readdata_pad_14.PULLUP = 1'b0;
    defparam readdata_pad_14.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_14.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_15 (.PACKAGE_PIN(readdata[15]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_15));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_15.PIN_TYPE = 6'b011001;
    defparam readdata_pad_15.PULLUP = 1'b0;
    defparam readdata_pad_15.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_15.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_16 (.PACKAGE_PIN(readdata[16]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_16));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_16.PIN_TYPE = 6'b011001;
    defparam readdata_pad_16.PULLUP = 1'b0;
    defparam readdata_pad_16.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_16.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_17 (.PACKAGE_PIN(readdata[17]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_17));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_17.PIN_TYPE = 6'b011001;
    defparam readdata_pad_17.PULLUP = 1'b0;
    defparam readdata_pad_17.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_17.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_18 (.PACKAGE_PIN(readdata[18]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_18));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_18.PIN_TYPE = 6'b011001;
    defparam readdata_pad_18.PULLUP = 1'b0;
    defparam readdata_pad_18.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_18.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_19 (.PACKAGE_PIN(readdata[19]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_19));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_19.PIN_TYPE = 6'b011001;
    defparam readdata_pad_19.PULLUP = 1'b0;
    defparam readdata_pad_19.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_19.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_20 (.PACKAGE_PIN(readdata[20]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_20));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_20.PIN_TYPE = 6'b011001;
    defparam readdata_pad_20.PULLUP = 1'b0;
    defparam readdata_pad_20.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_20.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_21 (.PACKAGE_PIN(readdata[21]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_21));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_21.PIN_TYPE = 6'b011001;
    defparam readdata_pad_21.PULLUP = 1'b0;
    defparam readdata_pad_21.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_21.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_22 (.PACKAGE_PIN(readdata[22]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_22));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_22.PIN_TYPE = 6'b011001;
    defparam readdata_pad_22.PULLUP = 1'b0;
    defparam readdata_pad_22.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_22.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_23 (.PACKAGE_PIN(readdata[23]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_23));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_23.PIN_TYPE = 6'b011001;
    defparam readdata_pad_23.PULLUP = 1'b0;
    defparam readdata_pad_23.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_23.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_24 (.PACKAGE_PIN(readdata[24]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_24));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_24.PIN_TYPE = 6'b011001;
    defparam readdata_pad_24.PULLUP = 1'b0;
    defparam readdata_pad_24.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_24.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_25 (.PACKAGE_PIN(readdata[25]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_25));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_25.PIN_TYPE = 6'b011001;
    defparam readdata_pad_25.PULLUP = 1'b0;
    defparam readdata_pad_25.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_25.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_26 (.PACKAGE_PIN(readdata[26]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_26));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_26.PIN_TYPE = 6'b011001;
    defparam readdata_pad_26.PULLUP = 1'b0;
    defparam readdata_pad_26.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_26.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_27 (.PACKAGE_PIN(readdata[27]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_27));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_27.PIN_TYPE = 6'b011001;
    defparam readdata_pad_27.PULLUP = 1'b0;
    defparam readdata_pad_27.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_27.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_28 (.PACKAGE_PIN(readdata[28]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_28));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_28.PIN_TYPE = 6'b011001;
    defparam readdata_pad_28.PULLUP = 1'b0;
    defparam readdata_pad_28.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_28.IO_STANDARD = "SB_LVCMOS";
    SB_IO readdata_pad_29 (.PACKAGE_PIN(readdata[29]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(readdata_c_29));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam readdata_pad_29.PIN_TYPE = 6'b011001;
    defparam readdata_pad_29.PULLUP = 1'b0;
    defparam readdata_pad_29.NEG_TRIGGER = 1'b0;
    defparam readdata_pad_29.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i7356_4_lut (.I0(ootx_payloads_1_181), .I1(data), .I2(n884), 
            .I3(lighthouse[0]), .O(n11466));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7356_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7357_4_lut (.I0(ootx_payloads_1_182), .I1(data), .I2(n886), 
            .I3(lighthouse[0]), .O(n11467));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7357_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i19_4_lut (.I0(counter_from_last_rise[31]), .I1(n6334), .I2(n2282), 
            .I3(n2), .O(n23397));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i19_4_lut_adj_886 (.I0(counter_from_last_rise[30]), .I1(n6335), 
            .I2(n2282), .I3(n2), .O(n23407));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i19_4_lut_adj_886.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_887 (.I0(counter_from_last_rise[29]), .I1(n6336), 
            .I2(n2282), .I3(n2), .O(n8_adj_2274));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_887.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_888 (.I0(counter_from_last_rise[28]), .I1(n6337), 
            .I2(n2282), .I3(n2), .O(n8_adj_2273));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_888.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_889 (.I0(counter_from_last_rise[27]), .I1(n6338), 
            .I2(n2282), .I3(n2), .O(n8_adj_2269));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_889.LUT_INIT = 16'h0aca;
    SB_LUT4 i7358_4_lut (.I0(ootx_payloads_1_183), .I1(data), .I2(n888), 
            .I3(lighthouse[0]), .O(n11468));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7358_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22_4_lut_adj_890 (.I0(counter_from_last_rise[26]), .I1(n6339), 
            .I2(n2282), .I3(n2), .O(n8_adj_2268));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_890.LUT_INIT = 16'h0aca;
    SB_LUT4 i7359_4_lut (.I0(ootx_payloads_1_184), .I1(data), .I2(n890), 
            .I3(lighthouse[0]), .O(n11469));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7359_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22_4_lut_adj_891 (.I0(counter_from_last_rise[25]), .I1(n6340), 
            .I2(n2282), .I3(n2), .O(n8_adj_2264));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_891.LUT_INIT = 16'h0aca;
    SB_LUT4 i7360_4_lut (.I0(ootx_payloads_1_185), .I1(data), .I2(n892), 
            .I3(lighthouse[0]), .O(n11470));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7360_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22_4_lut_adj_892 (.I0(counter_from_last_rise[24]), .I1(n6341), 
            .I2(n2282), .I3(n2), .O(n8_adj_2263));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_892.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_893 (.I0(counter_from_last_rise[23]), .I1(n6342), 
            .I2(n2282), .I3(n2), .O(n8_adj_2262));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_893.LUT_INIT = 16'h0aca;
    SB_LUT4 i7361_4_lut (.I0(ootx_payloads_1_186), .I1(data), .I2(n894), 
            .I3(lighthouse[0]), .O(n11471));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7361_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22_4_lut_adj_894 (.I0(counter_from_last_rise[22]), .I1(n6343), 
            .I2(n2282), .I3(n2), .O(n8_adj_2261));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_894.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_895 (.I0(counter_from_last_rise[21]), .I1(n6344), 
            .I2(n2282), .I3(n2), .O(n8_adj_2260));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_895.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_896 (.I0(counter_from_last_rise[20]), .I1(n6345), 
            .I2(n2282), .I3(n2), .O(n8_adj_2259));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_896.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_897 (.I0(counter_from_last_rise[19]), .I1(n6346), 
            .I2(n2282), .I3(n2), .O(n8_adj_2258));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_897.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_557_i9_3_lut (.I0(n4551[88]), .I1(n4551[104]), .I2(address_c_0), 
            .I3(GND_net), .O(n4157));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i9_4_lut (.I0(n25768), .I1(n4157), .I2(address_c_2), 
            .I3(address_c_1), .O(n3730));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_898 (.I0(counter_from_last_rise[18]), .I1(n6347), 
            .I2(n2282), .I3(n2), .O(n8_adj_2255));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_898.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_899 (.I0(counter_from_last_rise[17]), .I1(n6348), 
            .I2(n2282), .I3(n2), .O(n8_adj_2254));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_899.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_900 (.I0(counter_from_last_rise[16]), .I1(n6349), 
            .I2(n2282), .I3(n2), .O(n8_adj_2253));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_900.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_901 (.I0(counter_from_last_rise[15]), .I1(n6350), 
            .I2(n2282), .I3(n2), .O(n8_adj_2266));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_901.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_902 (.I0(counter_from_last_rise[14]), .I1(n6351), 
            .I2(n2282), .I3(n2), .O(n8_adj_2288));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_902.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_903 (.I0(counter_from_last_rise[13]), .I1(n6352), 
            .I2(n2282), .I3(n2), .O(n8_adj_2287));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_903.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_904 (.I0(counter_from_last_rise[12]), .I1(n6353), 
            .I2(n2282), .I3(n2), .O(n8_adj_2285));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_904.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_556_i10_3_lut (.I0(n4551[209]), .I1(n4551[225]), .I2(address_c_0), 
            .I3(GND_net), .O(n4139));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_567_i10_4_lut (.I0(n4139), .I1(n4551[241]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4302));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_905 (.I0(counter_from_last_rise[11]), .I1(n6354), 
            .I2(n2282), .I3(n2), .O(n8_adj_2282));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_905.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_553_i10_3_lut (.I0(n4551[137]), .I1(n4551[153]), .I2(address_c_0), 
            .I3(GND_net), .O(n4096));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_4_lut_adj_906 (.I0(counter_from_last_rise[10]), .I1(n6355), 
            .I2(n2282), .I3(n2), .O(n8_adj_2275));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_906.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_907 (.I0(counter_from_last_rise[9]), .I1(n6356), 
            .I2(n2282), .I3(n2), .O(n8_adj_2265));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_907.LUT_INIT = 16'h0aca;
    SB_LUT4 i20243_4_lut (.I0(\ootx_crc32_o[0] [16]), .I1(n7584), .I2(n4568[32]), 
            .I3(address_c_1), .O(n24616));
    defparam i20243_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15518167_i1_3_lut (.I0(n25540), .I1(n25396), .I2(address_c_2), 
            .I3(GND_net), .O(n3733));
    defparam i15518167_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_4_lut_adj_908 (.I0(counter_from_last_rise[8]), .I1(n6357), 
            .I2(n2282), .I3(n2), .O(n8_adj_2251));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_908.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_4_lut_adj_909 (.I0(counter_from_last_rise[7]), .I1(n6358), 
            .I2(n2282), .I3(n2), .O(n8));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_909.LUT_INIT = 16'h0aca;
    SB_LUT4 i7362_4_lut (.I0(ootx_payloads_1_187), .I1(data), .I2(n896), 
            .I3(lighthouse[0]), .O(n11472));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7362_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7363_4_lut (.I0(ootx_payloads_1_188), .I1(data), .I2(n898), 
            .I3(lighthouse[0]), .O(n11473));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7363_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7364_4_lut (.I0(ootx_payloads_1_189), .I1(data), .I2(n900), 
            .I3(lighthouse[0]), .O(n11474));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7364_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7365_4_lut (.I0(ootx_payloads_1_190), .I1(data), .I2(n902), 
            .I3(lighthouse[0]), .O(n11475));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7365_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22_4_lut_adj_910 (.I0(counter_from_last_rise[6]), .I1(n6359), 
            .I2(n2282), .I3(n2), .O(n8_adj_2296));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_910.LUT_INIT = 16'h0aca;
    SB_LUT4 i7366_4_lut (.I0(ootx_payloads_1_191), .I1(data), .I2(n904), 
            .I3(lighthouse[0]), .O(n11476));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7366_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7367_4_lut (.I0(ootx_payloads_1_192), .I1(data), .I2(n906), 
            .I3(lighthouse[0]), .O(n11477));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7367_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7368_4_lut (.I0(ootx_payloads_1_193), .I1(data), .I2(n908), 
            .I3(lighthouse[0]), .O(n11478));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7368_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7369_4_lut (.I0(ootx_payloads_1_194), .I1(data), .I2(n910), 
            .I3(lighthouse[0]), .O(n11479));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7369_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7370_4_lut (.I0(ootx_payloads_1_195), .I1(data), .I2(n912), 
            .I3(lighthouse[0]), .O(n11480));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7370_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22_4_lut_adj_911 (.I0(counter_from_last_rise[4]), .I1(n6361), 
            .I2(n2282), .I3(n2), .O(n8_adj_2281));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_911.LUT_INIT = 16'h0aca;
    SB_LUT4 i7371_4_lut (.I0(ootx_payloads_1_196), .I1(data), .I2(n914), 
            .I3(lighthouse[0]), .O(n11481));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7371_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7372_4_lut (.I0(ootx_payloads_1_197), .I1(data), .I2(n916), 
            .I3(lighthouse[0]), .O(n11482));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7372_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7373_4_lut (.I0(ootx_payloads_1_198), .I1(data), .I2(n918), 
            .I3(lighthouse[0]), .O(n11483));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7373_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7374_4_lut (.I0(ootx_payloads_1_199), .I1(data), .I2(n920), 
            .I3(lighthouse[0]), .O(n11484));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7374_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7375_4_lut (.I0(ootx_payloads_1_200), .I1(data), .I2(n922), 
            .I3(lighthouse[0]), .O(n11485));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7375_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7376_4_lut (.I0(ootx_payloads_1_201), .I1(data), .I2(n924), 
            .I3(lighthouse[0]), .O(n11486));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7376_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7377_4_lut (.I0(ootx_payloads_1_202), .I1(data), .I2(n926), 
            .I3(lighthouse[0]), .O(n11487));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7377_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_556_i11_3_lut (.I0(n4551[210]), .I1(n4551[226]), .I2(address_c_0), 
            .I3(GND_net), .O(n4138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_567_i11_4_lut (.I0(n4138), .I1(n4551[242]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4301));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7378_4_lut (.I0(ootx_payloads_1_203), .I1(data), .I2(n928), 
            .I3(lighthouse[0]), .O(n11488));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7378_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7379_4_lut (.I0(ootx_payloads_1_204), .I1(data), .I2(n930), 
            .I3(lighthouse[0]), .O(n11489));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7379_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7380_4_lut (.I0(ootx_payloads_1_205), .I1(data), .I2(n932), 
            .I3(lighthouse[0]), .O(n11490));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7380_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_553_i11_3_lut (.I0(n4551[138]), .I1(n4551[154]), .I2(address_c_0), 
            .I3(GND_net), .O(n4095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_556_i12_3_lut (.I0(n4551[211]), .I1(n4551[227]), .I2(address_c_0), 
            .I3(GND_net), .O(n4137));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_567_i12_4_lut (.I0(n4137), .I1(n4551[243]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4300));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7381_4_lut (.I0(ootx_payloads_1_206), .I1(data), .I2(n934), 
            .I3(lighthouse[0]), .O(n11491));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7381_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7382_4_lut (.I0(ootx_payloads_1_207), .I1(data), .I2(n936), 
            .I3(lighthouse[0]), .O(n11492));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7382_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_553_i12_3_lut (.I0(n4551[139]), .I1(n4551[155]), .I2(address_c_0), 
            .I3(GND_net), .O(n4094));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7383_4_lut (.I0(ootx_payloads_1_208), .I1(data), .I2(n938), 
            .I3(lighthouse[0]), .O(n11493));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7383_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7384_4_lut (.I0(ootx_payloads_1_209), .I1(data), .I2(n940), 
            .I3(lighthouse[0]), .O(n11494));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7384_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7385_4_lut (.I0(ootx_payloads_1_210), .I1(data), .I2(n942), 
            .I3(lighthouse[0]), .O(n11495));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7385_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7386_4_lut (.I0(ootx_payloads_1_211), .I1(data), .I2(n944), 
            .I3(lighthouse[0]), .O(n11496));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7386_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7387_4_lut (.I0(ootx_payloads_1_212), .I1(data), .I2(n946), 
            .I3(lighthouse[0]), .O(n11497));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7387_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7388_4_lut (.I0(ootx_payloads_1_213), .I1(data), .I2(n948), 
            .I3(lighthouse[0]), .O(n11498));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7388_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7389_4_lut (.I0(ootx_payloads_1_214), .I1(data), .I2(n950), 
            .I3(lighthouse[0]), .O(n11499));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7389_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7390_4_lut (.I0(ootx_payloads_1_215), .I1(data), .I2(n952), 
            .I3(lighthouse[0]), .O(n11500));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7390_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7391_4_lut (.I0(ootx_payloads_1_216), .I1(data), .I2(n954), 
            .I3(lighthouse[0]), .O(n11501));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7391_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7392_4_lut (.I0(ootx_payloads_1_217), .I1(data), .I2(n956), 
            .I3(lighthouse[0]), .O(n11502));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7392_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7393_4_lut (.I0(ootx_payloads_1_218), .I1(data), .I2(n958), 
            .I3(lighthouse[0]), .O(n11503));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7393_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i12_4_lut_adj_912 (.I0(data_counters_1_7), .I1(n361), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_912.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_913 (.I0(data_counters_1_6), .I1(n362), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_913.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_914 (.I0(data_counters_1_5), .I1(n363), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_914.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut (.I0(data_counters_1_4), .I1(n364), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_915 (.I0(data_counters_1_3), .I1(n365), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23071));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_915.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_916 (.I0(data_counters_1_2), .I1(n366), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23069));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_916.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_917 (.I0(data_counters_1_1), .I1(n367), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23067));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_917.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_918 (.I0(data_counters_1_0), .I1(n368), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23065));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_918.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_919 (.I0(data_counters_0_30), .I1(n338), .I2(n19), 
            .I3(n1), .O(n23063));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_919.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_920 (.I0(data_counters_0_29), .I1(n339), .I2(n19), 
            .I3(n1), .O(n23061));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_920.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_921 (.I0(data_counters_0_28), .I1(n340), .I2(n19), 
            .I3(n1), .O(n23059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_921.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_922 (.I0(data_counters_0_27), .I1(n341), .I2(n19), 
            .I3(n1), .O(n23057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_922.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_923 (.I0(data_counters_0_26), .I1(n342), .I2(n19), 
            .I3(n1), .O(n23055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_923.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_924 (.I0(data_counters_0_25), .I1(n343), .I2(n19), 
            .I3(n1), .O(n23053));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_924.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_925 (.I0(data_counters_0_24), .I1(n344), .I2(n19), 
            .I3(n1), .O(n23051));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_925.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_926 (.I0(data_counters_0_23), .I1(n345), .I2(n19), 
            .I3(n1), .O(n23049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_926.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_927 (.I0(data_counters_0_22), .I1(n346), .I2(n19), 
            .I3(n1), .O(n23047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_927.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_928 (.I0(data_counters_0_21), .I1(n347), .I2(n19), 
            .I3(n1), .O(n23045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_928.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_929 (.I0(data_counters_0_20), .I1(n348), .I2(n19), 
            .I3(n1), .O(n23043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_929.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_930 (.I0(data_counters_0_19), .I1(n349), .I2(n19), 
            .I3(n1), .O(n23041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_930.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_931 (.I0(data_counters_0_18), .I1(n350), .I2(n19), 
            .I3(n1), .O(n23039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_931.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_932 (.I0(data_counters_0_17), .I1(n351), .I2(n19), 
            .I3(n1), .O(n23037));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_932.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_933 (.I0(data_counters_0_16), .I1(n352), .I2(n19), 
            .I3(n1), .O(n23035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_933.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_934 (.I0(data_counters_0_15), .I1(n353), .I2(n19), 
            .I3(n1), .O(n23033));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_934.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_935 (.I0(data_counters_0_14), .I1(n354), .I2(n19), 
            .I3(n1), .O(n23031));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_935.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_936 (.I0(data_counters_0_13), .I1(n355), .I2(n19), 
            .I3(n1), .O(n23029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_936.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_937 (.I0(data_counters_0_12), .I1(n356), .I2(n19), 
            .I3(n1), .O(n23027));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_937.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_938 (.I0(data_counters_0_11), .I1(n357), .I2(n19), 
            .I3(n1), .O(n23025));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_938.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_939 (.I0(data_counters_0_10), .I1(n358), .I2(n19), 
            .I3(n1), .O(n23023));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_939.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_940 (.I0(data_counters_0_9), .I1(n359), .I2(n19), 
            .I3(n1), .O(n23021));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_940.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_941 (.I0(data_counters_0_8), .I1(n360), .I2(n19), 
            .I3(n1), .O(n23019));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_941.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_942 (.I0(data_counters_0_7), .I1(n361), .I2(n19), 
            .I3(n1), .O(n23017));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_942.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_943 (.I0(data_counters_0_6), .I1(n362), .I2(n19), 
            .I3(n1), .O(n23015));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_943.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_944 (.I0(data_counters_0_5), .I1(n363), .I2(n19), 
            .I3(n1), .O(n23013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_944.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_945 (.I0(data_counters_0_4), .I1(n364), .I2(n19), 
            .I3(n1), .O(n23011));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_945.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_946 (.I0(data_counters_0_3), .I1(n365), .I2(n19), 
            .I3(n1), .O(n23009));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_946.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_947 (.I0(data_counters_0_2), .I1(n366), .I2(n19), 
            .I3(n1), .O(n23007));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_947.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_948 (.I0(data_counters_0_1), .I1(n367), .I2(n19), 
            .I3(n1), .O(n23005));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_948.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_949 (.I0(data_counters_0_0), .I1(n368), .I2(n19), 
            .I3(n1), .O(n23003));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i11_4_lut_adj_949.LUT_INIT = 16'haca0;
    SB_LUT4 i46_4_lut (.I0(n23971), .I1(n28_adj_2276), .I2(ootx_payloads_N_1744[0]), 
            .I3(ootx_payloads_N_1698), .O(n25));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i46_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i45_4_lut (.I0(n13221), .I1(n25), .I2(ootx_payloads_N_1744[1]), 
            .I3(ootx_payloads_N_1744[0]), .O(n28_adj_2284));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i45_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 address_c_3_bdd_4_lut (.I0(address_c_3), .I1(n25822), .I2(n25348), 
            .I3(address_c_4), .O(n25885));
    defparam address_c_3_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25885_bdd_4_lut (.I0(n25885), .I1(n25306), .I2(n3728), .I3(address_c_4), 
            .O(n25888));
    defparam n25885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21098 (.I0(address_c_3), .I1(n25816), 
            .I2(n25354), .I3(address_c_4), .O(n25879));
    defparam address_c_3_bdd_4_lut_21098.LUT_INIT = 16'he4aa;
    SB_LUT4 n25879_bdd_4_lut (.I0(n25879), .I1(n25312), .I2(n3727), .I3(address_c_4), 
            .O(n25882));
    defparam n25879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21093 (.I0(address_c_3), .I1(n25810), 
            .I2(n25360), .I3(address_c_4), .O(n25873));
    defparam address_c_3_bdd_4_lut_21093.LUT_INIT = 16'he4aa;
    SB_LUT4 n25873_bdd_4_lut (.I0(n25873), .I1(n25318), .I2(n3726), .I3(address_c_4), 
            .O(n25876));
    defparam n25873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21088 (.I0(address_c_3), .I1(n25804), 
            .I2(n25366), .I3(address_c_4), .O(n25867));
    defparam address_c_3_bdd_4_lut_21088.LUT_INIT = 16'he4aa;
    SB_LUT4 n25867_bdd_4_lut (.I0(n25867), .I1(n25324), .I2(n3725), .I3(address_c_4), 
            .O(n25870));
    defparam n25867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21083 (.I0(address_c_3), .I1(n25798), 
            .I2(n25372), .I3(address_c_4), .O(n25861));
    defparam address_c_3_bdd_4_lut_21083.LUT_INIT = 16'he4aa;
    SB_LUT4 n25861_bdd_4_lut (.I0(n25861), .I1(n25330), .I2(n3724), .I3(address_c_4), 
            .O(n25864));
    defparam n25861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21078 (.I0(address_c_3), .I1(n25792), 
            .I2(n25378), .I3(address_c_4), .O(n25855));
    defparam address_c_3_bdd_4_lut_21078.LUT_INIT = 16'he4aa;
    SB_LUT4 n25855_bdd_4_lut (.I0(n25855), .I1(n25336), .I2(n3723), .I3(address_c_4), 
            .O(n25858));
    defparam n25855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21073 (.I0(address_c_3), .I1(n24832), 
            .I2(n24833), .I3(address_c_4), .O(n25849));
    defparam address_c_3_bdd_4_lut_21073.LUT_INIT = 16'he4aa;
    SB_LUT4 n25849_bdd_4_lut (.I0(n25849), .I1(n24654), .I2(n24653), .I3(address_c_4), 
            .O(n25852));
    defparam n25849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21068 (.I0(address_c_3), .I1(n24830), 
            .I2(n24831), .I3(address_c_4), .O(n25843));
    defparam address_c_3_bdd_4_lut_21068.LUT_INIT = 16'he4aa;
    SB_LUT4 n25843_bdd_4_lut (.I0(n25843), .I1(n24656), .I2(n24655), .I3(address_c_4), 
            .O(n25846));
    defparam n25843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_4_bdd_4_lut (.I0(address_c_4), .I1(n24825), .I2(n24826), 
            .I3(address_c_3), .O(n25837));
    defparam address_c_4_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25837_bdd_4_lut (.I0(n25837), .I1(n24658), .I2(n24657), .I3(address_c_3), 
            .O(n25840));
    defparam n25837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut (.I0(address_c_1), .I1(n4244), .I2(n4225), 
            .I3(address_c_2), .O(n25831));
    defparam address_c_1_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25831_bdd_4_lut (.I0(n25831), .I1(n3100), .I2(n24659), .I3(address_c_2), 
            .O(n24323));
    defparam n25831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21053 (.I0(address_c_1), .I1(n4243), .I2(n4224), 
            .I3(address_c_2), .O(n25825));
    defparam address_c_1_bdd_4_lut_21053.LUT_INIT = 16'he4aa;
    SB_LUT4 n25825_bdd_4_lut (.I0(n25825), .I1(n3099), .I2(n24660), .I3(address_c_2), 
            .O(n24326));
    defparam n25825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21048 (.I0(address_c_1), .I1(n4242), .I2(n4223), 
            .I3(address_c_2), .O(n25819));
    defparam address_c_1_bdd_4_lut_21048.LUT_INIT = 16'he4aa;
    SB_LUT4 n25819_bdd_4_lut (.I0(n25819), .I1(n3098), .I2(n24661), .I3(address_c_2), 
            .O(n25822));
    defparam n25819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21043 (.I0(address_c_1), .I1(n4241), .I2(n4222), 
            .I3(address_c_2), .O(n25813));
    defparam address_c_1_bdd_4_lut_21043.LUT_INIT = 16'he4aa;
    SB_LUT4 n25813_bdd_4_lut (.I0(n25813), .I1(n3097), .I2(n24662), .I3(address_c_2), 
            .O(n25816));
    defparam n25813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21038 (.I0(address_c_1), .I1(n4240), .I2(n4221), 
            .I3(address_c_2), .O(n25807));
    defparam address_c_1_bdd_4_lut_21038.LUT_INIT = 16'he4aa;
    SB_LUT4 n25807_bdd_4_lut (.I0(n25807), .I1(n3096), .I2(n24663), .I3(address_c_2), 
            .O(n25810));
    defparam n25807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21033 (.I0(address_c_1), .I1(n4239), .I2(n4220), 
            .I3(address_c_2), .O(n25801));
    defparam address_c_1_bdd_4_lut_21033.LUT_INIT = 16'he4aa;
    SB_LUT4 n25801_bdd_4_lut (.I0(n25801), .I1(n3095), .I2(n24664), .I3(address_c_2), 
            .O(n25804));
    defparam n25801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21028 (.I0(address_c_1), .I1(n4238), .I2(n4219), 
            .I3(address_c_2), .O(n25795));
    defparam address_c_1_bdd_4_lut_21028.LUT_INIT = 16'he4aa;
    SB_LUT4 n25795_bdd_4_lut (.I0(n25795), .I1(n3094), .I2(n24665), .I3(address_c_2), 
            .O(n25798));
    defparam n25795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21023 (.I0(address_c_1), .I1(n4237), .I2(n4218), 
            .I3(address_c_2), .O(n25789));
    defparam address_c_1_bdd_4_lut_21023.LUT_INIT = 16'he4aa;
    SB_LUT4 n25789_bdd_4_lut (.I0(n25789), .I1(n3093), .I2(n24666), .I3(address_c_2), 
            .O(n25792));
    defparam n25789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut (.I0(address_c_0), .I1(n4551[232]), .I2(n4551[248]), 
            .I3(address_c_1), .O(n25783));
    defparam address_c_0_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25783_bdd_4_lut (.I0(n25783), .I1(n4551[216]), .I2(n4551[200]), 
            .I3(address_c_1), .O(n24347));
    defparam n25783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_21013 (.I0(address_c_0), .I1(n4568[128]), 
            .I2(n4568[144]), .I3(address_c_1), .O(n25777));
    defparam address_c_0_bdd_4_lut_21013.LUT_INIT = 16'he4aa;
    SB_LUT4 n25777_bdd_4_lut (.I0(n25777), .I1(n4568[120]), .I2(n4568[112]), 
            .I3(address_c_1), .O(n24350));
    defparam n25777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_21008 (.I0(address_c_0), .I1(n4568[256]), 
            .I2(\ootx_crc32_o[1] [0]), .I3(address_c_1), .O(n25771));
    defparam address_c_0_bdd_4_lut_21008.LUT_INIT = 16'he4aa;
    SB_LUT4 n25771_bdd_4_lut (.I0(n25771), .I1(n4568[248]), .I2(n4568[232]), 
            .I3(address_c_1), .O(n25774));
    defparam n25771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_21003 (.I0(address_c_0), .I1(n4551[56]), 
            .I2(n4551[72]), .I3(address_c_1), .O(n25765));
    defparam address_c_0_bdd_4_lut_21003.LUT_INIT = 16'he4aa;
    SB_LUT4 n25765_bdd_4_lut (.I0(n25765), .I1(n4551[24]), .I2(n4551[8]), 
            .I3(address_c_1), .O(n25768));
    defparam n25765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20998 (.I0(address_c_0), .I1(n4551[57]), 
            .I2(n4551[73]), .I3(address_c_1), .O(n25759));
    defparam address_c_0_bdd_4_lut_20998.LUT_INIT = 16'he4aa;
    SB_LUT4 n25759_bdd_4_lut (.I0(n25759), .I1(n4551[25]), .I2(n4551[9]), 
            .I3(address_c_1), .O(n25762));
    defparam n25759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20993 (.I0(address_c_0), .I1(n4551[58]), 
            .I2(n4551[74]), .I3(address_c_1), .O(n25753));
    defparam address_c_0_bdd_4_lut_20993.LUT_INIT = 16'he4aa;
    SB_LUT4 n25753_bdd_4_lut (.I0(n25753), .I1(n4551[26]), .I2(n4551[10]), 
            .I3(address_c_1), .O(n25756));
    defparam n25753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20988 (.I0(address_c_0), .I1(n4551[59]), 
            .I2(n4551[75]), .I3(address_c_1), .O(n25747));
    defparam address_c_0_bdd_4_lut_20988.LUT_INIT = 16'he4aa;
    SB_LUT4 n25747_bdd_4_lut (.I0(n25747), .I1(n4551[27]), .I2(n4551[11]), 
            .I3(address_c_1), .O(n25750));
    defparam n25747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20983 (.I0(address_c_0), .I1(n4551[60]), 
            .I2(n4551[76]), .I3(address_c_1), .O(n25741));
    defparam address_c_0_bdd_4_lut_20983.LUT_INIT = 16'he4aa;
    SB_LUT4 n25741_bdd_4_lut (.I0(n25741), .I1(n4551[28]), .I2(n4551[12]), 
            .I3(address_c_1), .O(n25744));
    defparam n25741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20978 (.I0(address_c_0), .I1(n4551[61]), 
            .I2(n4551[77]), .I3(address_c_1), .O(n25735));
    defparam address_c_0_bdd_4_lut_20978.LUT_INIT = 16'he4aa;
    SB_LUT4 n25735_bdd_4_lut (.I0(n25735), .I1(n4551[29]), .I2(n4551[13]), 
            .I3(address_c_1), .O(n25738));
    defparam n25735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20973 (.I0(address_c_0), .I1(n4551[62]), 
            .I2(n4551[78]), .I3(address_c_1), .O(n25729));
    defparam address_c_0_bdd_4_lut_20973.LUT_INIT = 16'he4aa;
    SB_LUT4 n25729_bdd_4_lut (.I0(n25729), .I1(n4551[30]), .I2(n4551[14]), 
            .I3(address_c_1), .O(n25732));
    defparam n25729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20968 (.I0(address_c_0), .I1(n4551[63]), 
            .I2(n4551[79]), .I3(address_c_1), .O(n25723));
    defparam address_c_0_bdd_4_lut_20968.LUT_INIT = 16'he4aa;
    SB_LUT4 n25723_bdd_4_lut (.I0(n25723), .I1(n4551[31]), .I2(n4551[15]), 
            .I3(address_c_1), .O(n25726));
    defparam n25723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20963 (.I0(address_c_0), .I1(n4551[233]), 
            .I2(n4551[249]), .I3(address_c_1), .O(n25717));
    defparam address_c_0_bdd_4_lut_20963.LUT_INIT = 16'he4aa;
    SB_LUT4 n25717_bdd_4_lut (.I0(n25717), .I1(n4551[217]), .I2(n4551[201]), 
            .I3(address_c_1), .O(n24386));
    defparam n25717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20958 (.I0(address_c_0), .I1(n4551[234]), 
            .I2(n4551[250]), .I3(address_c_1), .O(n25711));
    defparam address_c_0_bdd_4_lut_20958.LUT_INIT = 16'he4aa;
    SB_LUT4 n25711_bdd_4_lut (.I0(n25711), .I1(n4551[218]), .I2(n4551[202]), 
            .I3(address_c_1), .O(n24389));
    defparam n25711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20953 (.I0(address_c_0), .I1(n4551[235]), 
            .I2(n4551[251]), .I3(address_c_1), .O(n25705));
    defparam address_c_0_bdd_4_lut_20953.LUT_INIT = 16'he4aa;
    SB_LUT4 n25705_bdd_4_lut (.I0(n25705), .I1(n4551[219]), .I2(n4551[203]), 
            .I3(address_c_1), .O(n24392));
    defparam n25705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20948 (.I0(address_c_0), .I1(n4551[236]), 
            .I2(n4551[252]), .I3(address_c_1), .O(n25699));
    defparam address_c_0_bdd_4_lut_20948.LUT_INIT = 16'he4aa;
    SB_LUT4 n25699_bdd_4_lut (.I0(n25699), .I1(n4551[220]), .I2(n4551[204]), 
            .I3(address_c_1), .O(n24398));
    defparam n25699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20943 (.I0(address_c_0), .I1(n4551[237]), 
            .I2(n4551[253]), .I3(address_c_1), .O(n25693));
    defparam address_c_0_bdd_4_lut_20943.LUT_INIT = 16'he4aa;
    SB_LUT4 n25693_bdd_4_lut (.I0(n25693), .I1(n4551[221]), .I2(n4551[205]), 
            .I3(address_c_1), .O(n24401));
    defparam n25693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20938 (.I0(address_c_0), .I1(n4551[238]), 
            .I2(n4551[254]), .I3(address_c_1), .O(n25687));
    defparam address_c_0_bdd_4_lut_20938.LUT_INIT = 16'he4aa;
    SB_LUT4 n25687_bdd_4_lut (.I0(n25687), .I1(n4551[222]), .I2(n4551[206]), 
            .I3(address_c_1), .O(n24404));
    defparam n25687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20933 (.I0(address_c_0), .I1(n4551[239]), 
            .I2(n4551[255]), .I3(address_c_1), .O(n25681));
    defparam address_c_0_bdd_4_lut_20933.LUT_INIT = 16'he4aa;
    SB_LUT4 n25681_bdd_4_lut (.I0(n25681), .I1(n4551[223]), .I2(n4551[207]), 
            .I3(address_c_1), .O(n24407));
    defparam n25681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20928 (.I0(address_c_0), .I1(n4568[129]), 
            .I2(n4568[145]), .I3(address_c_1), .O(n25675));
    defparam address_c_0_bdd_4_lut_20928.LUT_INIT = 16'he4aa;
    SB_LUT4 n25675_bdd_4_lut (.I0(n25675), .I1(n4568[121]), .I2(n4568[113]), 
            .I3(address_c_1), .O(n24410));
    defparam n25675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20923 (.I0(address_c_0), .I1(n4568[130]), 
            .I2(n4568[146]), .I3(address_c_1), .O(n25669));
    defparam address_c_0_bdd_4_lut_20923.LUT_INIT = 16'he4aa;
    SB_LUT4 n25669_bdd_4_lut (.I0(n25669), .I1(n4568[122]), .I2(n4568[114]), 
            .I3(address_c_1), .O(n24413));
    defparam n25669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20918 (.I0(address_c_0), .I1(n4568[131]), 
            .I2(n4568[147]), .I3(address_c_1), .O(n25663));
    defparam address_c_0_bdd_4_lut_20918.LUT_INIT = 16'he4aa;
    SB_LUT4 n25663_bdd_4_lut (.I0(n25663), .I1(n4568[123]), .I2(n4568[115]), 
            .I3(address_c_1), .O(n24416));
    defparam n25663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20913 (.I0(address_c_0), .I1(n4568[132]), 
            .I2(n4568[148]), .I3(address_c_1), .O(n25657));
    defparam address_c_0_bdd_4_lut_20913.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut (.I0(n28_adj_2284), .I1(lighthouse[0]), .I2(new_data), 
            .I3(GND_net), .O(n29));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n25657_bdd_4_lut (.I0(n25657), .I1(n4568[124]), .I2(n4568[116]), 
            .I3(address_c_1), .O(n24422));
    defparam n25657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20908 (.I0(address_c_0), .I1(n4568[133]), 
            .I2(n4568[149]), .I3(address_c_1), .O(n25651));
    defparam address_c_0_bdd_4_lut_20908.LUT_INIT = 16'he4aa;
    SB_LUT4 n25651_bdd_4_lut (.I0(n25651), .I1(n4568[125]), .I2(n4568[117]), 
            .I3(address_c_1), .O(n24425));
    defparam n25651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20903 (.I0(address_c_0), .I1(n4568[134]), 
            .I2(n4568[150]), .I3(address_c_1), .O(n25645));
    defparam address_c_0_bdd_4_lut_20903.LUT_INIT = 16'he4aa;
    SB_LUT4 n25645_bdd_4_lut (.I0(n25645), .I1(n4568[126]), .I2(n4568[118]), 
            .I3(address_c_1), .O(n24428));
    defparam n25645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20898 (.I0(address_c_0), .I1(n4568[135]), 
            .I2(n4568[151]), .I3(address_c_1), .O(n25639));
    defparam address_c_0_bdd_4_lut_20898.LUT_INIT = 16'he4aa;
    SB_LUT4 n25639_bdd_4_lut (.I0(n25639), .I1(n4568[127]), .I2(n4568[119]), 
            .I3(address_c_1), .O(n24431));
    defparam n25639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20893 (.I0(address_c_0), .I1(n4568[257]), 
            .I2(\ootx_crc32_o[1] [1]), .I3(address_c_1), .O(n25633));
    defparam address_c_0_bdd_4_lut_20893.LUT_INIT = 16'he4aa;
    SB_LUT4 n25633_bdd_4_lut (.I0(n25633), .I1(n4568[249]), .I2(n4568[233]), 
            .I3(address_c_1), .O(n25636));
    defparam n25633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20888 (.I0(address_c_0), .I1(n4568[258]), 
            .I2(\ootx_crc32_o[1] [2]), .I3(address_c_1), .O(n25627));
    defparam address_c_0_bdd_4_lut_20888.LUT_INIT = 16'he4aa;
    SB_LUT4 n25627_bdd_4_lut (.I0(n25627), .I1(n4568[250]), .I2(n4568[234]), 
            .I3(address_c_1), .O(n25630));
    defparam n25627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20883 (.I0(address_c_0), .I1(n4568[259]), 
            .I2(\ootx_crc32_o[1] [3]), .I3(address_c_1), .O(n25621));
    defparam address_c_0_bdd_4_lut_20883.LUT_INIT = 16'he4aa;
    SB_LUT4 n25621_bdd_4_lut (.I0(n25621), .I1(n4568[251]), .I2(n4568[235]), 
            .I3(address_c_1), .O(n25624));
    defparam n25621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut (.I0(n4702), .I1(n4568[169]), .I2(n4568[193]), 
            .I3(n4700), .O(n25615));
    defparam n4702_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25615_bdd_4_lut (.I0(n25615), .I1(n4079), .I2(n24627), .I3(n4700), 
            .O(n24179));
    defparam n25615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20878 (.I0(address_c_0), .I1(n4568[260]), 
            .I2(\ootx_crc32_o[1] [4]), .I3(address_c_1), .O(n25609));
    defparam address_c_0_bdd_4_lut_20878.LUT_INIT = 16'he4aa;
    SB_LUT4 n25609_bdd_4_lut (.I0(n25609), .I1(n4568[252]), .I2(n4568[236]), 
            .I3(address_c_1), .O(n25612));
    defparam n25609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20868 (.I0(address_c_0), .I1(n4568[261]), 
            .I2(\ootx_crc32_o[1] [5]), .I3(address_c_1), .O(n25603));
    defparam address_c_0_bdd_4_lut_20868.LUT_INIT = 16'he4aa;
    SB_LUT4 n25603_bdd_4_lut (.I0(n25603), .I1(n4568[253]), .I2(n4568[237]), 
            .I3(address_c_1), .O(n25606));
    defparam n25603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20873 (.I0(n4702), .I1(n4568[168]), .I2(n4568[192]), 
            .I3(n4700), .O(n25597));
    defparam n4702_bdd_4_lut_20873.LUT_INIT = 16'he4aa;
    SB_LUT4 n25597_bdd_4_lut (.I0(n25597), .I1(n4080), .I2(n24628), .I3(n4700), 
            .O(n24182));
    defparam n25597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20863 (.I0(address_c_0), .I1(n4568[262]), 
            .I2(\ootx_crc32_o[1] [6]), .I3(address_c_1), .O(n25591));
    defparam address_c_0_bdd_4_lut_20863.LUT_INIT = 16'he4aa;
    SB_LUT4 n25591_bdd_4_lut (.I0(n25591), .I1(n4568[254]), .I2(n4568[238]), 
            .I3(address_c_1), .O(n25594));
    defparam n25591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20853 (.I0(address_c_0), .I1(n4568[263]), 
            .I2(\ootx_crc32_o[1] [7]), .I3(address_c_1), .O(n25585));
    defparam address_c_0_bdd_4_lut_20853.LUT_INIT = 16'he4aa;
    SB_LUT4 n25585_bdd_4_lut (.I0(n25585), .I1(n4568[255]), .I2(n4568[239]), 
            .I3(address_c_1), .O(n25588));
    defparam n25585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20858 (.I0(n4702), .I1(n4568[167]), .I2(n4568[191]), 
            .I3(n4700), .O(n25579));
    defparam n4702_bdd_4_lut_20858.LUT_INIT = 16'he4aa;
    SB_LUT4 n25579_bdd_4_lut (.I0(n25579), .I1(n4081), .I2(n24431), .I3(n4700), 
            .O(n24185));
    defparam n25579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_21063 (.I0(address_c_3), .I1(n24800), 
            .I2(n24801), .I3(address_c_4), .O(n25573));
    defparam address_c_3_bdd_4_lut_21063.LUT_INIT = 16'he4aa;
    SB_LUT4 n25573_bdd_4_lut (.I0(n25573), .I1(n24725), .I2(n24724), .I3(address_c_4), 
            .O(n25576));
    defparam n25573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20838 (.I0(address_c_3), .I1(n24798), 
            .I2(n24799), .I3(address_c_4), .O(n25567));
    defparam address_c_3_bdd_4_lut_20838.LUT_INIT = 16'he4aa;
    SB_LUT4 n25567_bdd_4_lut (.I0(n25567), .I1(n24727), .I2(n24726), .I3(address_c_4), 
            .O(n25570));
    defparam n25567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20833 (.I0(address_c_3), .I1(n25456), 
            .I2(n25402), .I3(address_c_4), .O(n25561));
    defparam address_c_3_bdd_4_lut_20833.LUT_INIT = 16'he4aa;
    SB_LUT4 n25561_bdd_4_lut (.I0(n25561), .I1(n25390), .I2(n25462), .I3(address_c_4), 
            .O(n25564));
    defparam n25561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_4_bdd_4_lut_21058 (.I0(address_c_4), .I1(n24796), 
            .I2(n24797), .I3(address_c_3), .O(n25555));
    defparam address_c_4_bdd_4_lut_21058.LUT_INIT = 16'he4aa;
    SB_LUT4 n25555_bdd_4_lut (.I0(n25555), .I1(n24729), .I2(n24728), .I3(address_c_3), 
            .O(n25558));
    defparam n25555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i20475_4_lut (.I0(\ootx_states[1] [0]), .I1(n29), .I2(lighthouse[0]), 
            .I3(n23947), .O(n20_adj_2252));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i20475_4_lut.LUT_INIT = 16'h2232;
    SB_LUT4 address_c_4_bdd_4_lut_20823 (.I0(address_c_4), .I1(n24794), 
            .I2(n24795), .I3(address_c_3), .O(n25549));
    defparam address_c_4_bdd_4_lut_20823.LUT_INIT = 16'he4aa;
    SB_LUT4 n25549_bdd_4_lut (.I0(n25549), .I1(n24731), .I2(n24730), .I3(address_c_3), 
            .O(n25552));
    defparam n25549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut (.I0(n4673), .I1(n4551[161]), .I2(n4551[185]), 
            .I3(n4671), .O(n25543));
    defparam n4673_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25543_bdd_4_lut (.I0(n25543), .I1(n4104), .I2(n24386), .I3(n4671), 
            .O(n24152));
    defparam n25543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20848 (.I0(address_c_0), .I1(n4551[53]), 
            .I2(n4551[69]), .I3(address_c_1), .O(n25537));
    defparam address_c_0_bdd_4_lut_20848.LUT_INIT = 16'he4aa;
    SB_LUT4 n25537_bdd_4_lut (.I0(n25537), .I1(n4551[21]), .I2(n4551[5]), 
            .I3(address_c_1), .O(n25540));
    defparam n25537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20843 (.I0(n4702), .I1(n4568[166]), .I2(n4568[190]), 
            .I3(n4700), .O(n25531));
    defparam n4702_bdd_4_lut_20843.LUT_INIT = 16'he4aa;
    SB_LUT4 n25531_bdd_4_lut (.I0(n25531), .I1(n4082), .I2(n24428), .I3(n4700), 
            .O(n24188));
    defparam n25531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_21018 (.I0(address_c_1), .I1(n24147), 
            .I2(n24148), .I3(address_c_2), .O(n25525));
    defparam address_c_1_bdd_4_lut_21018.LUT_INIT = 16'he4aa;
    SB_LUT4 n25525_bdd_4_lut (.I0(n25525), .I1(n24514), .I2(n24513), .I3(address_c_2), 
            .O(n3734));
    defparam n25525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20799 (.I0(address_c_1), .I1(n24282), 
            .I2(n24283), .I3(address_c_2), .O(n25519));
    defparam address_c_1_bdd_4_lut_20799.LUT_INIT = 16'he4aa;
    SB_LUT4 n25519_bdd_4_lut (.I0(n25519), .I1(n24508), .I2(n24507), .I3(address_c_2), 
            .O(n3732));
    defparam n25519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20804 (.I0(n4702), .I1(n4568[165]), .I2(n4568[189]), 
            .I3(n4700), .O(n25513));
    defparam n4702_bdd_4_lut_20804.LUT_INIT = 16'he4aa;
    SB_LUT4 n25513_bdd_4_lut (.I0(n25513), .I1(n4083), .I2(n24425), .I3(n4700), 
            .O(n24191));
    defparam n25513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20794 (.I0(address_c_1), .I1(n24306), 
            .I2(n24307), .I3(address_c_2), .O(n25507));
    defparam address_c_1_bdd_4_lut_20794.LUT_INIT = 16'he4aa;
    SB_LUT4 n25507_bdd_4_lut (.I0(n25507), .I1(n24505), .I2(n24504), .I3(address_c_2), 
            .O(n3731));
    defparam n25507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20784 (.I0(address_c_1), .I1(n24309), 
            .I2(n24310), .I3(address_c_2), .O(n25501));
    defparam address_c_1_bdd_4_lut_20784.LUT_INIT = 16'he4aa;
    SB_LUT4 n25501_bdd_4_lut (.I0(n25501), .I1(n24502), .I2(n24501), .I3(address_c_2), 
            .O(n3805));
    defparam n25501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20779 (.I0(address_c_1), .I1(n24312), 
            .I2(n24313), .I3(address_c_2), .O(n25495));
    defparam address_c_1_bdd_4_lut_20779.LUT_INIT = 16'he4aa;
    SB_LUT4 n25495_bdd_4_lut (.I0(n25495), .I1(n24499), .I2(n24498), .I3(address_c_2), 
            .O(n3804));
    defparam n25495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20774 (.I0(address_c_1), .I1(n24315), 
            .I2(n24316), .I3(address_c_2), .O(n25489));
    defparam address_c_1_bdd_4_lut_20774.LUT_INIT = 16'he4aa;
    SB_LUT4 n25489_bdd_4_lut (.I0(n25489), .I1(n24496), .I2(n24495), .I3(address_c_2), 
            .O(n3803));
    defparam n25489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20769 (.I0(address_c_1), .I1(n24363), 
            .I2(n24364), .I3(address_c_2), .O(n25483));
    defparam address_c_1_bdd_4_lut_20769.LUT_INIT = 16'he4aa;
    SB_LUT4 n25483_bdd_4_lut (.I0(n25483), .I1(n24493), .I2(n24492), .I3(address_c_2), 
            .O(n3802));
    defparam n25483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20764 (.I0(address_c_1), .I1(n24366), 
            .I2(n24367), .I3(address_c_2), .O(n25477));
    defparam address_c_1_bdd_4_lut_20764.LUT_INIT = 16'he4aa;
    SB_LUT4 n25477_bdd_4_lut (.I0(n25477), .I1(n24490), .I2(n24489), .I3(address_c_2), 
            .O(n3801));
    defparam n25477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20759 (.I0(address_c_1), .I1(n24393), 
            .I2(n24394), .I3(address_c_2), .O(n25471));
    defparam address_c_1_bdd_4_lut_20759.LUT_INIT = 16'he4aa;
    SB_LUT4 n25471_bdd_4_lut (.I0(n25471), .I1(n24487), .I2(n24486), .I3(address_c_2), 
            .O(n3800));
    defparam n25471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20754 (.I0(address_c_1), .I1(n24417), 
            .I2(n24418), .I3(address_c_2), .O(n25465));
    defparam address_c_1_bdd_4_lut_20754.LUT_INIT = 16'he4aa;
    SB_LUT4 n25465_bdd_4_lut (.I0(n25465), .I1(n24469), .I2(n24468), .I3(address_c_2), 
            .O(n3799));
    defparam n25465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20749 (.I0(address_c_1), .I1(n24519), 
            .I2(n24520), .I3(address_c_2), .O(n25459));
    defparam address_c_1_bdd_4_lut_20749.LUT_INIT = 16'he4aa;
    SB_LUT4 n25459_bdd_4_lut (.I0(n25459), .I1(n24466), .I2(n24465), .I3(address_c_2), 
            .O(n25462));
    defparam n25459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20744 (.I0(address_c_1), .I1(n24522), 
            .I2(n24523), .I3(address_c_2), .O(n25453));
    defparam address_c_1_bdd_4_lut_20744.LUT_INIT = 16'he4aa;
    SB_LUT4 n25453_bdd_4_lut (.I0(n25453), .I1(n24463), .I2(n24462), .I3(address_c_2), 
            .O(n25456));
    defparam n25453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sensor_select_1__bdd_4_lut (.I0(sensor_select[1]), .I1(n24525), 
            .I2(n24526), .I3(sensor_select[2]), .O(n25447));
    defparam sensor_select_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n25447_bdd_4_lut (.I0(n25447), .I1(n24460), .I2(n24459), .I3(sensor_select[2]), 
            .O(sensor_N_132));
    defparam n25447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20739 (.I0(address_c_1), .I1(n24528), 
            .I2(n24529), .I3(address_c_2), .O(n25441));
    defparam address_c_1_bdd_4_lut_20739.LUT_INIT = 16'he4aa;
    SB_LUT4 n25441_bdd_4_lut (.I0(n25441), .I1(n24457), .I2(n24456), .I3(address_c_2), 
            .O(n3737));
    defparam n25441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20730 (.I0(address_c_1), .I1(n24531), 
            .I2(n24532), .I3(address_c_2), .O(n25435));
    defparam address_c_1_bdd_4_lut_20730.LUT_INIT = 16'he4aa;
    SB_LUT4 n25435_bdd_4_lut (.I0(n25435), .I1(n24454), .I2(n24453), .I3(address_c_2), 
            .O(n3736));
    defparam n25435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_1_bdd_4_lut_20725 (.I0(address_c_1), .I1(n24534), 
            .I2(n24535), .I3(address_c_2), .O(n25429));
    defparam address_c_1_bdd_4_lut_20725.LUT_INIT = 16'he4aa;
    SB_LUT4 n25429_bdd_4_lut (.I0(n25429), .I1(n24517), .I2(n24516), .I3(address_c_2), 
            .O(n3735));
    defparam n25429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20789 (.I0(n4702), .I1(n4568[164]), .I2(n4568[188]), 
            .I3(n4700), .O(n25423));
    defparam n4702_bdd_4_lut_20789.LUT_INIT = 16'he4aa;
    SB_LUT4 n25423_bdd_4_lut (.I0(n25423), .I1(n4084), .I2(n24422), .I3(n4700), 
            .O(n24194));
    defparam n25423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20716 (.I0(n4702), .I1(n4568[163]), .I2(n4568[187]), 
            .I3(n4700), .O(n25417));
    defparam n4702_bdd_4_lut_20716.LUT_INIT = 16'he4aa;
    SB_LUT4 n25417_bdd_4_lut (.I0(n25417), .I1(n4085), .I2(n24416), .I3(n4700), 
            .O(n24197));
    defparam n25417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20711 (.I0(n4702), .I1(n4568[162]), .I2(n4568[186]), 
            .I3(n4700), .O(n25411));
    defparam n4702_bdd_4_lut_20711.LUT_INIT = 16'he4aa;
    SB_LUT4 n25411_bdd_4_lut (.I0(n25411), .I1(n4086), .I2(n24413), .I3(n4700), 
            .O(n24200));
    defparam n25411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20706 (.I0(n4702), .I1(n4568[161]), .I2(n4568[185]), 
            .I3(n4700), .O(n25405));
    defparam n4702_bdd_4_lut_20706.LUT_INIT = 16'he4aa;
    SB_LUT4 n25405_bdd_4_lut (.I0(n25405), .I1(n4087), .I2(n24410), .I3(n4700), 
            .O(n24203));
    defparam n25405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20701 (.I0(n4702), .I1(n4568[160]), .I2(n4568[184]), 
            .I3(n4700), .O(n25399));
    defparam n4702_bdd_4_lut_20701.LUT_INIT = 16'he4aa;
    SB_LUT4 n25399_bdd_4_lut (.I0(n25399), .I1(n4088), .I2(n24350), .I3(n4700), 
            .O(n25402));
    defparam n25399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_0_bdd_4_lut_20809 (.I0(address_c_0), .I1(n4551[117]), 
            .I2(n4551[125]), .I3(address_c_1), .O(n25393));
    defparam address_c_0_bdd_4_lut_20809.LUT_INIT = 16'he4aa;
    SB_LUT4 n25393_bdd_4_lut (.I0(n25393), .I1(n4551[101]), .I2(n4551[85]), 
            .I3(address_c_1), .O(n25396));
    defparam n25393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20814 (.I0(n4673), .I1(n4551[160]), .I2(n4551[184]), 
            .I3(n4671), .O(n25387));
    defparam n4673_bdd_4_lut_20814.LUT_INIT = 16'he4aa;
    SB_LUT4 n25387_bdd_4_lut (.I0(n25387), .I1(n4105), .I2(n24347), .I3(n4671), 
            .O(n25390));
    defparam n25387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20687 (.I0(n4673), .I1(n4551[162]), .I2(n4551[186]), 
            .I3(n4671), .O(n25381));
    defparam n4673_bdd_4_lut_20687.LUT_INIT = 16'he4aa;
    SB_LUT4 n25381_bdd_4_lut (.I0(n25381), .I1(n4103), .I2(n24389), .I3(n4671), 
            .O(n24209));
    defparam n25381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20696 (.I0(n4702), .I1(n4568[175]), .I2(n4568[199]), 
            .I3(n4700), .O(n25375));
    defparam n4702_bdd_4_lut_20696.LUT_INIT = 16'he4aa;
    SB_LUT4 n25375_bdd_4_lut (.I0(n25375), .I1(n4073), .I2(n24620), .I3(n4700), 
            .O(n25378));
    defparam n25375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20677 (.I0(n4702), .I1(n4568[174]), .I2(n4568[198]), 
            .I3(n4700), .O(n25369));
    defparam n4702_bdd_4_lut_20677.LUT_INIT = 16'he4aa;
    SB_LUT4 n25369_bdd_4_lut (.I0(n25369), .I1(n4074), .I2(n24622), .I3(n4700), 
            .O(n25372));
    defparam n25369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20672 (.I0(n4702), .I1(n4568[173]), .I2(n4568[197]), 
            .I3(n4700), .O(n25363));
    defparam n4702_bdd_4_lut_20672.LUT_INIT = 16'he4aa;
    SB_LUT4 n25363_bdd_4_lut (.I0(n25363), .I1(n4075), .I2(n24623), .I3(n4700), 
            .O(n25366));
    defparam n25363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20667 (.I0(n4702), .I1(n4568[172]), .I2(n4568[196]), 
            .I3(n4700), .O(n25357));
    defparam n4702_bdd_4_lut_20667.LUT_INIT = 16'he4aa;
    SB_LUT4 n25357_bdd_4_lut (.I0(n25357), .I1(n4076), .I2(n24624), .I3(n4700), 
            .O(n25360));
    defparam n25357_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20662 (.I0(n4702), .I1(n4568[171]), .I2(n4568[195]), 
            .I3(n4700), .O(n25351));
    defparam n4702_bdd_4_lut_20662.LUT_INIT = 16'he4aa;
    SB_LUT4 n25351_bdd_4_lut (.I0(n25351), .I1(n4077), .I2(n24625), .I3(n4700), 
            .O(n25354));
    defparam n25351_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4702_bdd_4_lut_20657 (.I0(n4702), .I1(n4568[170]), .I2(n4568[194]), 
            .I3(n4700), .O(n25345));
    defparam n4702_bdd_4_lut_20657.LUT_INIT = 16'he4aa;
    SB_LUT4 n25345_bdd_4_lut (.I0(n25345), .I1(n4078), .I2(n24626), .I3(n4700), 
            .O(n25348));
    defparam n25345_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20682 (.I0(n4673), .I1(n4551[163]), .I2(n4551[187]), 
            .I3(n4671), .O(n25339));
    defparam n4673_bdd_4_lut_20682.LUT_INIT = 16'he4aa;
    SB_LUT4 n25339_bdd_4_lut (.I0(n25339), .I1(n4102), .I2(n24392), .I3(n4671), 
            .O(n24212));
    defparam n25339_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20648 (.I0(n4673), .I1(n4551[175]), .I2(n4551[199]), 
            .I3(n4671), .O(n25333));
    defparam n4673_bdd_4_lut_20648.LUT_INIT = 16'he4aa;
    SB_LUT4 n25333_bdd_4_lut (.I0(n25333), .I1(n4090), .I2(n4296), .I3(n4671), 
            .O(n25336));
    defparam n25333_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20643 (.I0(n4673), .I1(n4551[174]), .I2(n4551[198]), 
            .I3(n4671), .O(n25327));
    defparam n4673_bdd_4_lut_20643.LUT_INIT = 16'he4aa;
    SB_LUT4 n25327_bdd_4_lut (.I0(n25327), .I1(n4091), .I2(n4297), .I3(n4671), 
            .O(n25330));
    defparam n25327_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20638 (.I0(n4673), .I1(n4551[173]), .I2(n4551[197]), 
            .I3(n4671), .O(n25321));
    defparam n4673_bdd_4_lut_20638.LUT_INIT = 16'he4aa;
    SB_LUT4 n25321_bdd_4_lut (.I0(n25321), .I1(n4092), .I2(n4298), .I3(n4671), 
            .O(n25324));
    defparam n25321_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n4673_bdd_4_lut_20633 (.I0(n4673), .I1(n4551[172]), .I2(n4551[196]), 
            .I3(n4671), .O(n25315));
    defparam n4673_bdd_4_lut_20633.LUT_INIT = 16'he4aa;
    SB_LUT4 n25315_bdd_4_lut (.I0(n25315), .I1(n4093), .I2(n4299), .I3(n4671), 
            .O(n25318));
    defparam n25315_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7394_4_lut (.I0(ootx_payloads_1_219), .I1(data), .I2(n960), 
            .I3(lighthouse[0]), .O(n11504));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7394_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7395_4_lut (.I0(ootx_payloads_1_220), .I1(data), .I2(n962), 
            .I3(lighthouse[0]), .O(n11505));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7395_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), .I2(address_c_3), 
            .I3(address_c_2), .O(n13397));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i20267_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[32]), .I3(address_c_2), .O(n24634));
    defparam i20267_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20279_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[36]), .I3(address_c_2), .O(n24730));
    defparam i20279_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20451_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[33]), .I3(address_c_2), .O(n24728));
    defparam i20451_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20453_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[39]), .I3(address_c_2), .O(n24726));
    defparam i20453_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20455_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[38]), .I3(address_c_2), .O(n24657));
    defparam i20455_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20256_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[37]), .I3(address_c_2), .O(n24724));
    defparam i20256_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20456_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[35]), .I3(address_c_2), .O(n24655));
    defparam i20456_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i20271_2_lut_3_lut_4_lut (.I0(address_c_0), .I1(address_c_1), 
            .I2(n4551[34]), .I3(address_c_2), .O(n24653));
    defparam i20271_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i7396_4_lut (.I0(ootx_payloads_1_221), .I1(data), .I2(n964), 
            .I3(lighthouse[0]), .O(n11506));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7396_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_950 (.I0(address_c_2), .I1(address_c_0), .I2(GND_net), 
            .I3(GND_net), .O(n7584));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h4444;
    SB_LUT4 i20396_2_lut (.I0(n4568[47]), .I1(address_c_4), .I2(GND_net), 
            .I3(GND_net), .O(n24815));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i20396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7397_4_lut (.I0(ootx_payloads_1_222), .I1(data), .I2(n966), 
            .I3(lighthouse[0]), .O(n11507));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7397_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7398_4_lut (.I0(ootx_payloads_1_223), .I1(data), .I2(n968), 
            .I3(lighthouse[0]), .O(n11508));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7398_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_557_i10_3_lut (.I0(n4551[89]), .I1(n4551[105]), .I2(address_c_0), 
            .I3(GND_net), .O(n4156));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_557_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_529_i10_4_lut (.I0(n25762), .I1(n4156), .I2(address_c_2), 
            .I3(address_c_1), .O(n3729));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_529_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7399_4_lut (.I0(ootx_payloads_1_224), .I1(data), .I2(n970), 
            .I3(lighthouse[0]), .O(n11509));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7399_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i9321_3_lut (.I0(n4551[47]), .I1(\ootx_crc32_o[0] [31]), .I2(address_c_4), 
            .I3(GND_net), .O(n13426));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i9321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20426_4_lut (.I0(n13426), .I1(n50_adj_2283), .I2(n24815), 
            .I3(address_c_1), .O(n24782));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20426_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14896_4_lut (.I0(n24782), .I1(n72), .I2(n24783), .I3(address_c_5), 
            .O(readdata_c_31));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14896_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i7400_4_lut (.I0(ootx_payloads_1_225), .I1(data), .I2(n972), 
            .I3(lighthouse[0]), .O(n11510));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7400_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7401_4_lut (.I0(ootx_payloads_1_226), .I1(data), .I2(n974), 
            .I3(lighthouse[0]), .O(n11511));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7401_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7402_4_lut (.I0(ootx_payloads_1_227), .I1(data), .I2(n976), 
            .I3(lighthouse[0]), .O(n11512));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7402_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7403_4_lut (.I0(ootx_payloads_1_228), .I1(data), .I2(n978), 
            .I3(lighthouse[0]), .O(n11513));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7403_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7404_4_lut (.I0(ootx_payloads_1_229), .I1(data), .I2(n980), 
            .I3(lighthouse[0]), .O(n11514));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7404_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7405_4_lut (.I0(ootx_payloads_1_230), .I1(data), .I2(n982), 
            .I3(lighthouse[0]), .O(n11515));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7405_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7406_4_lut (.I0(ootx_payloads_1_231), .I1(data), .I2(n984), 
            .I3(lighthouse[0]), .O(n11516));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7406_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7407_4_lut (.I0(ootx_payloads_1_232), .I1(data), .I2(n986), 
            .I3(lighthouse[0]), .O(n11517));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7407_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7408_4_lut (.I0(ootx_payloads_1_233), .I1(data), .I2(n988), 
            .I3(lighthouse[0]), .O(n11518));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7408_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7409_4_lut (.I0(ootx_payloads_1_234), .I1(data), .I2(n990), 
            .I3(lighthouse[0]), .O(n11519));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7409_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7410_4_lut (.I0(ootx_payloads_1_235), .I1(data), .I2(n992), 
            .I3(lighthouse[0]), .O(n11520));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7410_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7411_4_lut (.I0(ootx_payloads_1_236), .I1(data), .I2(n994), 
            .I3(lighthouse[0]), .O(n11521));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7411_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFFER sensor_select__0__i2 (.Q(sensor_select[1]), .C(clock_c), .E(n2208), 
            .D(writedata_c_1), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(103[11] 109[5])
    SB_DFFER sensor_select__0__i3 (.Q(sensor_select[2]), .C(clock_c), .E(n2208), 
            .D(writedata_c_2), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(103[11] 109[5])
    SB_LUT4 i7412_4_lut (.I0(ootx_payloads_1_237), .I1(data), .I2(n996), 
            .I3(lighthouse[0]), .O(n11522));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7412_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7413_4_lut (.I0(ootx_payloads_1_238), .I1(data), .I2(n998), 
            .I3(lighthouse[0]), .O(n11523));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7413_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7414_4_lut (.I0(ootx_payloads_1_239), .I1(data), .I2(n1000), 
            .I3(lighthouse[0]), .O(n11524));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7414_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7415_4_lut (.I0(ootx_payloads_1_240), .I1(data), .I2(n1002), 
            .I3(lighthouse[0]), .O(n11525));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7415_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7416_4_lut (.I0(ootx_payloads_1_241), .I1(data), .I2(n1004), 
            .I3(lighthouse[0]), .O(n11526));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7416_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7417_4_lut (.I0(ootx_payloads_1_242), .I1(data), .I2(n1006), 
            .I3(lighthouse[0]), .O(n11527));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7417_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7418_4_lut (.I0(ootx_payloads_1_243), .I1(data), .I2(n1008), 
            .I3(lighthouse[0]), .O(n11528));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7418_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7419_4_lut (.I0(ootx_payloads_1_244), .I1(data), .I2(n1010), 
            .I3(lighthouse[0]), .O(n11529));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7419_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7420_4_lut (.I0(ootx_payloads_1_245), .I1(data), .I2(n1012), 
            .I3(lighthouse[0]), .O(n11530));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7420_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7421_4_lut (.I0(ootx_payloads_1_246), .I1(data), .I2(n1014), 
            .I3(lighthouse[0]), .O(n11531));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7421_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7422_4_lut (.I0(ootx_payloads_1_247), .I1(data), .I2(n1016), 
            .I3(lighthouse[0]), .O(n11532));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7422_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7423_4_lut (.I0(ootx_payloads_1_248), .I1(data), .I2(n1018), 
            .I3(lighthouse[0]), .O(n11533));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7423_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7424_4_lut (.I0(ootx_payloads_1_249), .I1(data), .I2(n1020), 
            .I3(lighthouse[0]), .O(n11534));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7424_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7425_4_lut (.I0(ootx_payloads_1_250), .I1(data), .I2(n1022), 
            .I3(lighthouse[0]), .O(n11535));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7425_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7426_4_lut (.I0(ootx_payloads_1_251), .I1(data), .I2(n1024), 
            .I3(lighthouse[0]), .O(n11536));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7426_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7427_4_lut (.I0(ootx_payloads_1_252), .I1(data), .I2(n1026), 
            .I3(lighthouse[0]), .O(n11537));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7427_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7428_4_lut (.I0(ootx_payloads_1_253), .I1(data), .I2(n1028), 
            .I3(lighthouse[0]), .O(n11538));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7428_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7429_4_lut (.I0(ootx_payloads_1_254), .I1(data), .I2(n1030), 
            .I3(lighthouse[0]), .O(n11539));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7429_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7430_4_lut (.I0(ootx_payloads_1_255), .I1(data), .I2(n1032), 
            .I3(lighthouse[0]), .O(n11540));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7430_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7431_4_lut (.I0(ootx_payloads_1_256), .I1(data), .I2(n521), 
            .I3(lighthouse[0]), .O(n11541));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7431_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7432_4_lut (.I0(ootx_payloads_1_257), .I1(data), .I2(n523), 
            .I3(lighthouse[0]), .O(n11542));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7432_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7433_4_lut (.I0(ootx_payloads_1_258), .I1(data), .I2(n525), 
            .I3(lighthouse[0]), .O(n11543));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7433_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7434_4_lut (.I0(ootx_payloads_1_259), .I1(data), .I2(n527), 
            .I3(lighthouse[0]), .O(n11544));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7434_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7435_4_lut (.I0(ootx_payloads_1_260), .I1(data), .I2(n529), 
            .I3(lighthouse[0]), .O(n11545));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7435_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7436_4_lut (.I0(ootx_payloads_1_261), .I1(data), .I2(n531), 
            .I3(lighthouse[0]), .O(n11546));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7436_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7437_4_lut (.I0(ootx_payloads_1_262), .I1(data), .I2(n533), 
            .I3(lighthouse[0]), .O(n11547));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7437_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7438_4_lut (.I0(ootx_payloads_1_263), .I1(data), .I2(n535), 
            .I3(lighthouse[0]), .O(n11548));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i7438_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7439_4_lut (.I0(crc32s_1_0), .I1(data), .I2(n38), .I3(lighthouse[0]), 
            .O(n11549));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7439_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7440_4_lut (.I0(crc32s_1_1), .I1(data), .I2(n40), .I3(lighthouse[0]), 
            .O(n11550));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7440_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7441_4_lut (.I0(crc32s_1_2), .I1(data), .I2(n42), .I3(lighthouse[0]), 
            .O(n11551));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7441_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7442_4_lut (.I0(crc32s_1_3), .I1(data), .I2(n44), .I3(lighthouse[0]), 
            .O(n11552));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7442_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7443_4_lut (.I0(crc32s_1_4), .I1(data), .I2(n46), .I3(lighthouse[0]), 
            .O(n11553));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7443_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7444_4_lut (.I0(crc32s_1_5), .I1(data), .I2(n48), .I3(lighthouse[0]), 
            .O(n11554));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7444_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7445_4_lut (.I0(crc32s_1_6), .I1(data), .I2(n50), .I3(lighthouse[0]), 
            .O(n11555));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7445_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7446_4_lut (.I0(crc32s_1_7), .I1(data), .I2(n52), .I3(lighthouse[0]), 
            .O(n11556));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7446_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7447_4_lut (.I0(crc32s_1_8), .I1(data), .I2(n54_adj_2272), 
            .I3(lighthouse[0]), .O(n11557));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7447_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7448_4_lut (.I0(crc32s_1_9), .I1(data), .I2(n56), .I3(lighthouse[0]), 
            .O(n11558));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7448_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7449_4_lut (.I0(crc32s_1_10), .I1(data), .I2(n58), .I3(lighthouse[0]), 
            .O(n11559));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7449_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7450_4_lut (.I0(crc32s_1_11), .I1(data), .I2(n60), .I3(lighthouse[0]), 
            .O(n11560));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7450_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7451_4_lut (.I0(crc32s_1_12), .I1(data), .I2(n62), .I3(lighthouse[0]), 
            .O(n11561));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7451_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7452_4_lut (.I0(crc32s_1_13), .I1(data), .I2(n64), .I3(lighthouse[0]), 
            .O(n11562));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7452_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7453_4_lut (.I0(crc32s_1_14), .I1(data), .I2(n66), .I3(lighthouse[0]), 
            .O(n11563));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7453_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7454_4_lut (.I0(crc32s_1_15), .I1(data), .I2(n68), .I3(lighthouse[0]), 
            .O(n11564));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7454_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7455_4_lut (.I0(crc32s_1_16), .I1(data), .I2(n37_adj_2270), 
            .I3(lighthouse[0]), .O(n11565));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7455_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7456_4_lut (.I0(crc32s_1_17), .I1(data), .I2(n39), .I3(lighthouse[0]), 
            .O(n11566));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7456_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7457_4_lut (.I0(crc32s_1_18), .I1(data), .I2(n41), .I3(lighthouse[0]), 
            .O(n11567));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7457_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7458_4_lut (.I0(crc32s_1_19), .I1(data), .I2(n43), .I3(lighthouse[0]), 
            .O(n11568));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7458_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7459_4_lut (.I0(crc32s_1_20), .I1(data), .I2(n45_adj_2271), 
            .I3(lighthouse[0]), .O(n11569));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7459_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_951 (.I0(ootx_payloads_N_1744[0]), .I1(new_data), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(n35_adj_2257), .I1(n4), .I2(ootx_payloads_N_1698), 
            .I3(ootx_payloads_N_1744[1]), .O(n23947));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i2_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 n4673_bdd_4_lut_20628 (.I0(n4673), .I1(n4551[171]), .I2(n4551[195]), 
            .I3(n4671), .O(n25309));
    defparam n4673_bdd_4_lut_20628.LUT_INIT = 16'he4aa;
    SB_LUT4 i19393_2_lut (.I0(n13), .I1(lighthouse[0]), .I2(GND_net), 
            .I3(GND_net), .O(n24030));
    defparam i19393_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7460_4_lut (.I0(crc32s_1_21), .I1(data), .I2(n47), .I3(lighthouse[0]), 
            .O(n11570));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7460_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7461_4_lut (.I0(crc32s_1_22), .I1(data), .I2(n49), .I3(lighthouse[0]), 
            .O(n11571));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7461_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i20169_3_lut (.I0(lighthouse[0]), .I1(n23974), .I2(data), 
            .I3(GND_net), .O(n24540));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i20169_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i7462_4_lut (.I0(crc32s_1_23), .I1(data), .I2(n51), .I3(lighthouse[0]), 
            .O(n11572));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7462_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7463_4_lut (.I0(crc32s_1_24), .I1(data), .I2(n53), .I3(lighthouse[0]), 
            .O(n11573));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7463_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7464_4_lut (.I0(crc32s_1_25), .I1(data), .I2(n55), .I3(lighthouse[0]), 
            .O(n11574));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7464_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n24540), .I1(n24030), .I2(ootx_payloads_N_1744[1]), 
            .I3(n24018), .O(n33));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i53_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 n25309_bdd_4_lut (.I0(n25309), .I1(n4094), .I2(n4300), .I3(n4671), 
            .O(n25312));
    defparam n25309_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut (.I0(lighthouse[0]), .I1(n30_adj_2286), .I2(\ootx_states[0] [1]), 
            .I3(n23971), .O(n23972));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i3_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i7465_4_lut (.I0(crc32s_1_26), .I1(data), .I2(n57), .I3(lighthouse[0]), 
            .O(n11575));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7465_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut (.I0(new_data), .I1(n23972), .I2(ootx_payloads_N_1744[0]), 
            .I3(n33), .O(n37));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i1_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 n4673_bdd_4_lut_20623 (.I0(n4673), .I1(n4551[170]), .I2(n4551[194]), 
            .I3(n4671), .O(n25303));
    defparam n4673_bdd_4_lut_20623.LUT_INIT = 16'he4aa;
    SB_LUT4 i7466_4_lut (.I0(crc32s_1_27), .I1(data), .I2(n59), .I3(lighthouse[0]), 
            .O(n11576));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7466_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7467_4_lut (.I0(crc32s_1_28), .I1(data), .I2(n61), .I3(lighthouse[0]), 
            .O(n11577));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7467_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i20472_4_lut (.I0(\ootx_states[0] [0]), .I1(n37), .I2(lighthouse[0]), 
            .I3(n23947), .O(n25_adj_2299));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i20472_4_lut.LUT_INIT = 16'h2223;
    SB_LUT4 i7468_4_lut (.I0(crc32s_1_29), .I1(data), .I2(n63), .I3(lighthouse[0]), 
            .O(n11578));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7468_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n25303_bdd_4_lut (.I0(n25303), .I1(n4095), .I2(n4301), .I3(n4671), 
            .O(n25306));
    defparam n25303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7469_4_lut (.I0(crc32s_1_30), .I1(data), .I2(n65), .I3(lighthouse[0]), 
            .O(n11579));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7469_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7470_4_lut (.I0(crc32s_1_31), .I1(data), .I2(n67), .I3(lighthouse[0]), 
            .O(n11580));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7470_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i7471_4_lut (.I0(n3111), .I1(data), .I2(n38), .I3(lighthouse[0]), 
            .O(n11581));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7471_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7472_4_lut (.I0(n3110), .I1(data), .I2(n40), .I3(lighthouse[0]), 
            .O(n11582));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7472_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 n4673_bdd_4_lut_20618 (.I0(n4673), .I1(n4551[169]), .I2(n4551[193]), 
            .I3(n4671), .O(n25297));
    defparam n4673_bdd_4_lut_20618.LUT_INIT = 16'he4aa;
    SB_LUT4 i7473_4_lut (.I0(n3109), .I1(data), .I2(n42), .I3(lighthouse[0]), 
            .O(n11583));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7473_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7474_4_lut (.I0(n3108), .I1(data), .I2(n44), .I3(lighthouse[0]), 
            .O(n11584));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7474_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7475_4_lut (.I0(n3107), .I1(data), .I2(n46), .I3(lighthouse[0]), 
            .O(n11585));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7475_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 n25297_bdd_4_lut (.I0(n25297), .I1(n4096), .I2(n4302), .I3(n4671), 
            .O(n24233));
    defparam n25297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7476_4_lut (.I0(n3106), .I1(data), .I2(n48), .I3(lighthouse[0]), 
            .O(n11586));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7476_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7477_4_lut (.I0(n3105), .I1(data), .I2(n50), .I3(lighthouse[0]), 
            .O(n11587));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7477_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7478_4_lut (.I0(n3104), .I1(data), .I2(n52), .I3(lighthouse[0]), 
            .O(n11588));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7478_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7479_4_lut (.I0(n3103), .I1(data), .I2(n54_adj_2272), .I3(lighthouse[0]), 
            .O(n11589));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7479_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7480_4_lut (.I0(n3102), .I1(data), .I2(n56), .I3(lighthouse[0]), 
            .O(n11590));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7480_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7481_4_lut (.I0(n3101), .I1(data), .I2(n58), .I3(lighthouse[0]), 
            .O(n11591));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7481_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7482_4_lut (.I0(n3100_adj_2250), .I1(data), .I2(n60), .I3(lighthouse[0]), 
            .O(n11592));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7482_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7483_4_lut (.I0(n3099_adj_2249), .I1(data), .I2(n62), .I3(lighthouse[0]), 
            .O(n11593));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7483_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7484_4_lut (.I0(n3098_adj_2248), .I1(data), .I2(n64), .I3(lighthouse[0]), 
            .O(n11594));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7484_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7485_4_lut (.I0(n3097_adj_2247), .I1(data), .I2(n66), .I3(lighthouse[0]), 
            .O(n11595));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7485_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7486_4_lut (.I0(n3096_adj_2246), .I1(data), .I2(n68), .I3(lighthouse[0]), 
            .O(n11596));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7486_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i7487_4_lut (.I0(n3095_adj_2245), .I1(data), .I2(n37_adj_2270), 
            .I3(lighthouse[0]), .O(n11597));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7487_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i22_4_lut_adj_952 (.I0(counter_from_last_rise[3]), .I1(n6362), 
            .I2(reset_c), .I3(n2), .O(n8_adj_2277));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_952.LUT_INIT = 16'ha0ac;
    SB_LUT4 i7488_4_lut (.I0(n3094_adj_2244), .I1(data), .I2(n39), .I3(lighthouse[0]), 
            .O(n11598));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7488_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i22_4_lut_adj_953 (.I0(counter_from_last_rise[2]), .I1(n6363), 
            .I2(reset_c), .I3(n2), .O(n8_adj_2278));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_953.LUT_INIT = 16'ha0ac;
    SB_LUT4 i22_4_lut_adj_954 (.I0(counter_from_last_rise[1]), .I1(n6364), 
            .I2(reset_c), .I3(n2), .O(n8_adj_2279));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i22_4_lut_adj_954.LUT_INIT = 16'ha0ac;
    SB_LUT4 i1_4_lut_adj_955 (.I0(n35), .I1(payload_lengths_1_0), .I2(data), 
            .I3(n17), .O(n23641));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'h5044;
    SB_LUT4 i7489_4_lut (.I0(n3093_adj_2243), .I1(data), .I2(n41), .I3(lighthouse[0]), 
            .O(n11599));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7489_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i1_4_lut_adj_956 (.I0(n36), .I1(data), .I2(payload_lengths_0_0), 
            .I3(n19468), .O(n23639));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam i1_4_lut_adj_956.LUT_INIT = 16'h5044;
    SB_LUT4 i7490_4_lut (.I0(n3092), .I1(data), .I2(n43), .I3(lighthouse[0]), 
            .O(n11600));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7490_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12_4_lut_adj_957 (.I0(new_data), .I1(n24692), .I2(reset_c), 
            .I3(data_N_1808), .O(n23697));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i12_4_lut_adj_957.LUT_INIT = 16'haca0;
    SB_LUT4 i11_4_lut_adj_958 (.I0(bit_counters_1_30), .I1(n2852), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23391));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_958.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_959 (.I0(bit_counters_1_29), .I1(n2853), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23401));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_959.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_960 (.I0(n3091), .I1(data), .I2(lighthouse[0]), 
            .I3(n45_adj_2271), .O(n23001));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(50[9:13])
    defparam i11_4_lut_adj_960.LUT_INIT = 16'hacaa;
    SB_LUT4 i11_4_lut_adj_961 (.I0(bit_counters_1_28), .I1(n2854), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23411));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_961.LUT_INIT = 16'hca0a;
    SB_LUT4 i7492_4_lut (.I0(n3090), .I1(data), .I2(n47), .I3(lighthouse[0]), 
            .O(n11602));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7492_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i11_4_lut_adj_962 (.I0(bit_counters_1_27), .I1(n2855), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23417));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_962.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_963 (.I0(bit_counters_1_26), .I1(n2856), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23423));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_963.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_964 (.I0(n3089), .I1(data), .I2(lighthouse[0]), 
            .I3(n49), .O(n22997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(50[9:13])
    defparam i11_4_lut_adj_964.LUT_INIT = 16'hacaa;
    SB_LUT4 i12_4_lut_adj_965 (.I0(bit_counters_1_25), .I1(n2857), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23429));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_965.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_966 (.I0(bit_counters_1_24), .I1(n2858), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23435));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_966.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_967 (.I0(bit_counters_1_23), .I1(n2859), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23441));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_967.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_968 (.I0(bit_counters_1_22), .I1(n2860), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23447));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_968.LUT_INIT = 16'hca0a;
    SB_LUT4 i7494_4_lut (.I0(n3088), .I1(data), .I2(n51), .I3(lighthouse[0]), 
            .O(n11604));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7494_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12_4_lut_adj_969 (.I0(bit_counters_1_21), .I1(n2861), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23453));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_969.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_970 (.I0(bit_counters_1_20), .I1(n2862), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23459));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_970.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_971 (.I0(bit_counters_1_19), .I1(n2863), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23465));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_971.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_972 (.I0(bit_counters_1_18), .I1(n2864), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23471));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_972.LUT_INIT = 16'hca0a;
    SB_LUT4 i7495_4_lut (.I0(n3087), .I1(data), .I2(n53), .I3(lighthouse[0]), 
            .O(n11605));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7495_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 n4673_bdd_4_lut_20613 (.I0(n4673), .I1(n4551[168]), .I2(n4551[192]), 
            .I3(n4671), .O(n25291));
    defparam n4673_bdd_4_lut_20613.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_973 (.I0(bit_counters_1_17), .I1(n2865), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23545));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_973.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_974 (.I0(bit_counters_1_16), .I1(n2866), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23543));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_974.LUT_INIT = 16'hca0a;
    SB_LUT4 n25291_bdd_4_lut (.I0(n25291), .I1(n4097), .I2(n4303), .I3(n4671), 
            .O(n24236));
    defparam n25291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_975 (.I0(bit_counters_1_15), .I1(n2867), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23541));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_975.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_976 (.I0(bit_counters_1_14), .I1(n2868), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23539));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_976.LUT_INIT = 16'hca0a;
    SB_LUT4 i7496_4_lut (.I0(n3086), .I1(data), .I2(n55), .I3(lighthouse[0]), 
            .O(n11606));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7496_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12_4_lut_adj_977 (.I0(bit_counters_1_13), .I1(n2869), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23537));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_977.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_978 (.I0(bit_counters_1_12), .I1(n2870), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23535));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_978.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_979 (.I0(bit_counters_1_11), .I1(n2871), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23533));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_979.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_980 (.I0(bit_counters_1_10), .I1(n2872), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23531));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_980.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_981 (.I0(bit_counters_1_9), .I1(n2873), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23529));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_981.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_982 (.I0(bit_counters_1_8), .I1(n2874), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23527));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_982.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_983 (.I0(bit_counters_1_7), .I1(n2875), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23525));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_983.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_984 (.I0(bit_counters_1_6), .I1(n2876), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23523));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_984.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_985 (.I0(bit_counters_1_5), .I1(n2877), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23521));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_985.LUT_INIT = 16'hca0a;
    SB_LUT4 i7497_4_lut (.I0(n3085), .I1(data), .I2(n57), .I3(lighthouse[0]), 
            .O(n11607));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7497_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12_4_lut_adj_986 (.I0(bit_counters_1_4), .I1(n2878), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23519));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_986.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_987 (.I0(bit_counters_1_3), .I1(n2879), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23517));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_987.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_988 (.I0(bit_counters_1_2), .I1(n2880), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23515));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_988.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_989 (.I0(bit_counters_1_1), .I1(n2881), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23513));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_989.LUT_INIT = 16'hca0a;
    SB_LUT4 i7498_4_lut (.I0(n3084), .I1(data), .I2(n59), .I3(lighthouse[0]), 
            .O(n11608));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7498_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 n4673_bdd_4_lut_20608 (.I0(n4673), .I1(n4551[167]), .I2(n4551[191]), 
            .I3(n4671), .O(n25285));
    defparam n4673_bdd_4_lut_20608.LUT_INIT = 16'he4aa;
    SB_LUT4 i7499_4_lut (.I0(n3083), .I1(data), .I2(n61), .I3(lighthouse[0]), 
            .O(n11609));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7499_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12_4_lut_adj_990 (.I0(bit_counters_1_0), .I1(n2882), .I2(n9797), 
            .I3(n1_adj_2256), .O(n23511));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_990.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_991 (.I0(bit_counters_0_30), .I1(n2852), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23389));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_991.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_992 (.I0(bit_counters_0_29), .I1(n2853), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23399));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_992.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_993 (.I0(bit_counters_0_28), .I1(n2854), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23409));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_993.LUT_INIT = 16'hca0a;
    SB_LUT4 i7500_4_lut (.I0(n3082), .I1(data), .I2(n63), .I3(lighthouse[0]), 
            .O(n11610));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7500_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i11_4_lut_adj_994 (.I0(bit_counters_0_27), .I1(n2855), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23415));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_994.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_995 (.I0(bit_counters_0_26), .I1(n2856), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23421));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i11_4_lut_adj_995.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_996 (.I0(bit_counters_0_25), .I1(n2857), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23427));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_996.LUT_INIT = 16'hca0a;
    SB_LUT4 n25285_bdd_4_lut (.I0(n25285), .I1(n4098), .I2(n24407), .I3(n4671), 
            .O(n24239));
    defparam n25285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_997 (.I0(bit_counters_0_24), .I1(n2858), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23433));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_997.LUT_INIT = 16'hca0a;
    SB_LUT4 i7501_4_lut (.I0(n3081), .I1(data), .I2(n65), .I3(lighthouse[0]), 
            .O(n11611));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7501_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12_4_lut_adj_998 (.I0(bit_counters_0_23), .I1(n2859), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23439));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_998.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_999 (.I0(bit_counters_0_22), .I1(n2860), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23445));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_999.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1000 (.I0(bit_counters_0_21), .I1(n2861), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23451));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1000.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1001 (.I0(bit_counters_0_20), .I1(n2862), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23457));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1001.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1002 (.I0(bit_counters_0_19), .I1(n2863), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23463));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1002.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1003 (.I0(bit_counters_0_18), .I1(n2864), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23469));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1003.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1004 (.I0(bit_counters_0_17), .I1(n2865), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23509));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1004.LUT_INIT = 16'hca0a;
    SB_LUT4 i7502_4_lut (.I0(n3080), .I1(data), .I2(n67), .I3(lighthouse[0]), 
            .O(n11612));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    defparam i7502_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 n4673_bdd_4_lut_20603 (.I0(n4673), .I1(n4551[166]), .I2(n4551[190]), 
            .I3(n4671), .O(n25279));
    defparam n4673_bdd_4_lut_20603.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_1005 (.I0(bit_counters_0_16), .I1(n2866), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23507));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1005.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1006 (.I0(bit_counters_0_15), .I1(n2867), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23505));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1006.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1007 (.I0(bit_counters_0_14), .I1(n2868), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23503));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1007.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1008 (.I0(bit_counters_0_13), .I1(n2869), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23501));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1008.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1009 (.I0(bit_counters_0_12), .I1(n2870), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23499));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1009.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1010 (.I0(bit_counters_0_11), .I1(n2871), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23497));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1010.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1011 (.I0(bit_counters_0_10), .I1(n2872), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23495));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1011.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1012 (.I0(bit_counters_0_9), .I1(n2873), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23493));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1012.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1013 (.I0(bit_counters_0_8), .I1(n2874), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23491));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1013.LUT_INIT = 16'hca0a;
    SB_LUT4 n25279_bdd_4_lut (.I0(n25279), .I1(n4099), .I2(n24404), .I3(n4671), 
            .O(n24242));
    defparam n25279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1014 (.I0(bit_counters_0_7), .I1(n2875), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23489));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1014.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1015 (.I0(bit_counters_0_6), .I1(n2876), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23487));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1015.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1016 (.I0(bit_counters_0_5), .I1(n2877), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23485));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1016.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1017 (.I0(bit_counters_0_4), .I1(n2878), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23483));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1017.LUT_INIT = 16'hca0a;
    SB_LUT4 n4673_bdd_4_lut_20598 (.I0(n4673), .I1(n4551[165]), .I2(n4551[189]), 
            .I3(n4671), .O(n25273));
    defparam n4673_bdd_4_lut_20598.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_1018 (.I0(bit_counters_0_3), .I1(n2879), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23481));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1018.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1019 (.I0(bit_counters_0_2), .I1(n2880), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23479));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1019.LUT_INIT = 16'hca0a;
    SB_LUT4 n25273_bdd_4_lut (.I0(n25273), .I1(n4100), .I2(n24401), .I3(n4671), 
            .O(n24245));
    defparam n25273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1020 (.I0(bit_counters_0_1), .I1(n2881), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23477));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1020.LUT_INIT = 16'hca0a;
    SB_LUT4 n4673_bdd_4_lut_20593 (.I0(n4673), .I1(n4551[164]), .I2(n4551[188]), 
            .I3(n4671), .O(n25267));
    defparam n4673_bdd_4_lut_20593.LUT_INIT = 16'he4aa;
    SB_LUT4 n25267_bdd_4_lut (.I0(n25267), .I1(n4101), .I2(n24398), .I3(n4671), 
            .O(n24248));
    defparam n25267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1021 (.I0(bit_counters_0_0), .I1(n2882), .I2(n9771), 
            .I3(n1_adj_2267), .O(n23475));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    defparam i12_4_lut_adj_1021.LUT_INIT = 16'hca0a;
    SB_LUT4 i12_4_lut_adj_1022 (.I0(data_counters_1_30), .I1(n338), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1022.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1023 (.I0(data_counters_1_29), .I1(n339), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1023.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1024 (.I0(data_counters_1_28), .I1(n340), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23121));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1024.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1025 (.I0(data_counters_1_27), .I1(n341), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1025.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1026 (.I0(data_counters_1_26), .I1(n342), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1026.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1027 (.I0(data_counters_1_25), .I1(n343), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23115));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1027.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1028 (.I0(data_counters_1_24), .I1(n344), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1028.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1029 (.I0(data_counters_1_23), .I1(n345), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1029.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1030 (.I0(data_counters_1_22), .I1(n346), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1030.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1031 (.I0(data_counters_1_21), .I1(n347), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1031.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1032 (.I0(data_counters_1_20), .I1(n348), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1032.LUT_INIT = 16'haca0;
    SB_LUT4 i12_4_lut_adj_1033 (.I0(data_counters_1_19), .I1(n349), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1033.LUT_INIT = 16'haca0;
    SB_LUT4 mux_556_i13_3_lut (.I0(n4551[212]), .I1(n4551[228]), .I2(address_c_0), 
            .I3(GND_net), .O(n4136));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut (.I0(writedata_c_21), .I1(writedata_c_28), .I2(writedata_c_26), 
            .I3(writedata_c_19), .O(n44_adj_2298));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(writedata_c_30), .I1(writedata_c_14), .I2(writedata_c_22), 
            .I3(writedata_c_3), .O(n43_adj_2297));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(writedata_c_13), .I1(writedata_c_8), .I2(writedata_c_29), 
            .I3(writedata_c_5), .O(n49_adj_2289));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(writedata_c_4), .I1(writedata_c_7), .I2(writedata_c_10), 
            .I3(writedata_c_9), .O(n48_adj_2295));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(writedata_c_12), .I1(writedata_c_24), .I2(writedata_c_16), 
            .I3(writedata_c_18), .O(n46_adj_2292));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1034 (.I0(writedata_c_11), .I1(writedata_c_17), 
            .I2(writedata_c_15), .I3(writedata_c_20), .O(n47_adj_2293));
    defparam i19_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(writedata_c_23), .I1(writedata_c_27), .I2(writedata_c_25), 
            .I3(writedata_c_6), .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_adj_2293), .I2(n46_adj_2292), 
            .I3(n48_adj_2295), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_3_lut (.I0(n49_adj_2289), .I1(n43_adj_2297), .I2(n44_adj_2298), 
            .I3(GND_net), .O(n53_adj_2294));
    defparam i25_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(writedata_c_31), .I1(address_c_4), .I2(n53_adj_2294), 
            .I3(n54), .O(n7));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'h2223;
    SB_LUT4 i3_4_lut_adj_1036 (.I0(address_c_0), .I1(address_c_1), .I2(address_c_3), 
            .I3(address_c_2), .O(n9));
    defparam i3_4_lut_adj_1036.LUT_INIT = 16'h0001;
    SB_LUT4 i5_4_lut (.I0(n9), .I1(n7), .I2(write_c), .I3(address_c_5), 
            .O(n2208));
    defparam i5_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 mux_567_i13_4_lut (.I0(n4136), .I1(n4551[244]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4299));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_4_lut_adj_1037 (.I0(data_counters_1_18), .I1(n350), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1037.LUT_INIT = 16'haca0;
    SB_LUT4 mux_553_i13_3_lut (.I0(n4551[140]), .I1(n4551[156]), .I2(address_c_0), 
            .I3(GND_net), .O(n4093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1038 (.I0(data_counters_1_17), .I1(n351), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1038.LUT_INIT = 16'haca0;
    SB_LUT4 mux_556_i14_3_lut (.I0(n4551[213]), .I1(n4551[229]), .I2(address_c_0), 
            .I3(GND_net), .O(n4135));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1039 (.I0(data_counters_1_16), .I1(n352), .I2(n20_adj_2290), 
            .I3(n1_adj_2291), .O(n23097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i12_4_lut_adj_1039.LUT_INIT = 16'haca0;
    SB_LUT4 mux_567_i14_4_lut (.I0(n4135), .I1(n4551[245]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4298));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_553_i14_3_lut (.I0(n4551[141]), .I1(n4551[157]), .I2(address_c_0), 
            .I3(GND_net), .O(n4092));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_556_i15_3_lut (.I0(n4551[214]), .I1(n4551[230]), .I2(address_c_0), 
            .I3(GND_net), .O(n4134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_567_i15_4_lut (.I0(n4134), .I1(n4551[246]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4297));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_553_i15_3_lut (.I0(n4551[142]), .I1(n4551[158]), .I2(address_c_0), 
            .I3(GND_net), .O(n4091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_556_i16_3_lut (.I0(n4551[215]), .I1(n4551[231]), .I2(address_c_0), 
            .I3(GND_net), .O(n4133));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_556_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_567_i16_4_lut (.I0(n4133), .I1(n4551[247]), .I2(address_c_1), 
            .I3(address_c_0), .O(n4296));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_567_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_553_i16_3_lut (.I0(n4551[143]), .I1(n4551[159]), .I2(address_c_0), 
            .I3(GND_net), .O(n4090));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_553_i4_3_lut (.I0(n4551[131]), .I1(n4551[147]), .I2(address_c_0), 
            .I3(GND_net), .O(n4102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20368_4_lut (.I0(n4568[138]), .I1(address_c_1), .I2(n4568[154]), 
            .I3(address_c_0), .O(n24626));
    defparam i20368_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i11_3_lut (.I0(n4568[210]), .I1(n4568[226]), .I2(address_c_0), 
            .I3(GND_net), .O(n4078));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20369_4_lut (.I0(n4568[139]), .I1(address_c_1), .I2(n4568[155]), 
            .I3(address_c_0), .O(n24625));
    defparam i20369_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i12_3_lut (.I0(n4568[211]), .I1(n4568[227]), .I2(address_c_0), 
            .I3(GND_net), .O(n4077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20402_4_lut (.I0(\ootx_crc32_o[0] [29]), .I1(n8917), .I2(n4568[45]), 
            .I3(address_c_1), .O(n24765));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20402_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_541_i30_4_lut (.I0(n4551[45]), .I1(n24765), .I2(address_c_4), 
            .I3(n13397), .O(n3913));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_541_i30_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i14894_4_lut (.I0(n3913), .I1(n72), .I2(n24780), .I3(address_c_5), 
            .O(readdata_c_29));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14894_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i20370_4_lut (.I0(n4568[140]), .I1(address_c_1), .I2(n4568[156]), 
            .I3(address_c_0), .O(n24624));
    defparam i20370_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20394_2_lut (.I0(n4568[44]), .I1(address_c_4), .I2(GND_net), 
            .I3(GND_net), .O(n24812));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i20394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_552_i13_3_lut (.I0(n4568[212]), .I1(n4568[228]), .I2(address_c_0), 
            .I3(GND_net), .O(n4076));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9297_3_lut (.I0(n4551[44]), .I1(\ootx_crc32_o[0] [28]), .I2(address_c_4), 
            .I3(GND_net), .O(n13402));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i9297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20429_4_lut (.I0(n13402), .I1(n50_adj_2283), .I2(n24812), 
            .I3(address_c_1), .O(n24778));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20429_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14893_4_lut (.I0(n24778), .I1(n72), .I2(n24779), .I3(address_c_5), 
            .O(readdata_c_28));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14893_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i20371_4_lut (.I0(n4568[141]), .I1(address_c_1), .I2(n4568[157]), 
            .I3(address_c_0), .O(n24623));
    defparam i20371_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20401_4_lut (.I0(\ootx_crc32_o[0] [27]), .I1(n8917), .I2(n4568[43]), 
            .I3(address_c_1), .O(n24763));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20401_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i14_3_lut (.I0(n4568[213]), .I1(n4568[229]), .I2(address_c_0), 
            .I3(GND_net), .O(n4075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_541_i28_4_lut (.I0(n4551[43]), .I1(n24763), .I2(address_c_4), 
            .I3(n13397), .O(n3915));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_541_i28_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i14892_4_lut (.I0(n3915), .I1(n72), .I2(n24777), .I3(address_c_5), 
            .O(readdata_c_27));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14892_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i20246_4_lut (.I0(n4568[142]), .I1(address_c_1), .I2(n4568[158]), 
            .I3(address_c_0), .O(n24622));
    defparam i20246_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20403_4_lut (.I0(\ootx_crc32_o[0] [26]), .I1(n8917), .I2(n4568[42]), 
            .I3(address_c_1), .O(n24761));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20403_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i15_3_lut (.I0(n4568[214]), .I1(n4568[230]), .I2(address_c_0), 
            .I3(GND_net), .O(n4074));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20245_4_lut (.I0(n4568[143]), .I1(address_c_1), .I2(n4568[159]), 
            .I3(address_c_0), .O(n24620));
    defparam i20245_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_541_i27_4_lut (.I0(n4551[42]), .I1(n24761), .I2(address_c_4), 
            .I3(n13397), .O(n3916));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_541_i27_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 address_c_3_bdd_4_lut_20828 (.I0(address_c_3), .I1(n3805), .I2(n24203), 
            .I3(address_c_4), .O(n25261));
    defparam address_c_3_bdd_4_lut_20828.LUT_INIT = 16'he4aa;
    SB_LUT4 n25261_bdd_4_lut (.I0(n25261), .I1(n24152), .I2(n3737), .I3(address_c_4), 
            .O(n25264));
    defparam n25261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20584 (.I0(address_c_3), .I1(n3804), .I2(n24200), 
            .I3(address_c_4), .O(n25255));
    defparam address_c_3_bdd_4_lut_20584.LUT_INIT = 16'he4aa;
    SB_LUT4 n25255_bdd_4_lut (.I0(n25255), .I1(n24209), .I2(n3736), .I3(address_c_4), 
            .O(n25258));
    defparam n25255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20579 (.I0(address_c_3), .I1(n3803), .I2(n24197), 
            .I3(address_c_4), .O(n25249));
    defparam address_c_3_bdd_4_lut_20579.LUT_INIT = 16'he4aa;
    SB_LUT4 n25249_bdd_4_lut (.I0(n25249), .I1(n24212), .I2(n3735), .I3(address_c_4), 
            .O(n25252));
    defparam n25249_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20574 (.I0(address_c_3), .I1(n3802), .I2(n24194), 
            .I3(address_c_4), .O(n25243));
    defparam address_c_3_bdd_4_lut_20574.LUT_INIT = 16'he4aa;
    SB_LUT4 n25243_bdd_4_lut (.I0(n25243), .I1(n24248), .I2(n3734), .I3(address_c_4), 
            .O(n25246));
    defparam n25243_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20569 (.I0(address_c_3), .I1(n3801), .I2(n24191), 
            .I3(address_c_4), .O(n25237));
    defparam address_c_3_bdd_4_lut_20569.LUT_INIT = 16'he4aa;
    SB_LUT4 n25237_bdd_4_lut (.I0(n25237), .I1(n24245), .I2(n3733), .I3(address_c_4), 
            .O(n25240));
    defparam n25237_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20564 (.I0(address_c_3), .I1(n24616), 
            .I2(n24617), .I3(address_c_4), .O(n25231));
    defparam address_c_3_bdd_4_lut_20564.LUT_INIT = 16'he4aa;
    SB_LUT4 n25231_bdd_4_lut (.I0(n25231), .I1(n24635), .I2(n24634), .I3(address_c_4), 
            .O(n25234));
    defparam n25231_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20559 (.I0(address_c_3), .I1(n3800), .I2(n24188), 
            .I3(address_c_4), .O(n25225));
    defparam address_c_3_bdd_4_lut_20559.LUT_INIT = 16'he4aa;
    SB_LUT4 n25225_bdd_4_lut (.I0(n25225), .I1(n24242), .I2(n3732), .I3(address_c_4), 
            .O(n25228));
    defparam n25225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20554 (.I0(address_c_3), .I1(n3799), .I2(n24185), 
            .I3(address_c_4), .O(n25213));
    defparam address_c_3_bdd_4_lut_20554.LUT_INIT = 16'he4aa;
    SB_LUT4 n25213_bdd_4_lut (.I0(n25213), .I1(n24239), .I2(n3731), .I3(address_c_4), 
            .O(n25216));
    defparam n25213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 address_c_3_bdd_4_lut_20545 (.I0(address_c_3), .I1(n24323), 
            .I2(n24182), .I3(address_c_4), .O(n25207));
    defparam address_c_3_bdd_4_lut_20545.LUT_INIT = 16'he4aa;
    SB_LUT4 n25207_bdd_4_lut (.I0(n25207), .I1(n24236), .I2(n3730), .I3(address_c_4), 
            .O(n25210));
    defparam n25207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14891_4_lut (.I0(n3916), .I1(n72), .I2(n24776), .I3(address_c_5), 
            .O(readdata_c_26));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14891_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i20405_4_lut (.I0(\ootx_crc32_o[0] [25]), .I1(n8917), .I2(n4568[41]), 
            .I3(address_c_1), .O(n24759));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20405_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i16_3_lut (.I0(n4568[215]), .I1(n4568[231]), .I2(address_c_0), 
            .I3(GND_net), .O(n4073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_541_i26_4_lut (.I0(n4551[41]), .I1(n24759), .I2(address_c_4), 
            .I3(n13397), .O(n3917));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_541_i26_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i14890_4_lut (.I0(n3917), .I1(n72), .I2(n24775), .I3(address_c_5), 
            .O(readdata_c_25));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14890_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i20395_2_lut (.I0(n4568[40]), .I1(address_c_4), .I2(GND_net), 
            .I3(GND_net), .O(n24814));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i20395_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9309_3_lut (.I0(n4551[40]), .I1(\ootx_crc32_o[0] [24]), .I2(address_c_4), 
            .I3(GND_net), .O(n13414));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i9309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20433_4_lut (.I0(n13414), .I1(n50_adj_2283), .I2(n24814), 
            .I3(address_c_1), .O(n24773));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20433_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14889_4_lut (.I0(n24773), .I1(n72), .I2(n24774), .I3(address_c_5), 
            .O(readdata_c_24));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14889_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i14888_4_lut (.I0(n25570), .I1(n72), .I2(n24772), .I3(address_c_5), 
            .O(readdata_c_23));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14888_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1040 (.I0(n72), .I1(n25840), .I2(n24639), .I3(address_c_5), 
            .O(readdata_c_22));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'h5044;
    SB_LUT4 i14887_4_lut (.I0(n25576), .I1(n72), .I2(n24771), .I3(address_c_5), 
            .O(readdata_c_21));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14887_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1041 (.I0(n72), .I1(n25552), .I2(n24642), .I3(address_c_5), 
            .O(readdata_c_20));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'h5044;
    SB_LUT4 mux_553_i3_3_lut (.I0(n4551[130]), .I1(n4551[146]), .I2(address_c_0), 
            .I3(GND_net), .O(n4103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14886_4_lut (.I0(n25846), .I1(n72), .I2(n24770), .I3(address_c_5), 
            .O(readdata_c_19));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14886_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14885_4_lut (.I0(n25852), .I1(n72), .I2(n24769), .I3(address_c_5), 
            .O(readdata_c_18));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14885_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_553_i1_3_lut (.I0(n4551[128]), .I1(n4551[144]), .I2(address_c_0), 
            .I3(GND_net), .O(n4105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_552_i1_3_lut (.I0(n4568[200]), .I1(n4568[216]), .I2(address_c_0), 
            .I3(GND_net), .O(n4088));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(n72), .I1(n25558), .I2(n24643), .I3(address_c_5), 
            .O(readdata_c_17));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'h5044;
    SB_LUT4 address_c_3_bdd_4_lut_20540 (.I0(address_c_3), .I1(n24326), 
            .I2(n24179), .I3(address_c_4), .O(n25201));
    defparam address_c_3_bdd_4_lut_20540.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_552_i2_3_lut (.I0(n4568[201]), .I1(n4568[217]), .I2(address_c_0), 
            .I3(GND_net), .O(n4087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_552_i3_3_lut (.I0(n4568[202]), .I1(n4568[218]), .I2(address_c_0), 
            .I3(GND_net), .O(n4086));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14884_4_lut (.I0(n25234), .I1(n72), .I2(n24768), .I3(address_c_5), 
            .O(readdata_c_16));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14884_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_527_i16_4_lut (.I0(n4568[247]), .I1(\ootx_crc32_o[1] [15]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3689));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i16_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i14883_4_lut (.I0(n25858), .I1(n72), .I2(n3689), .I3(address_c_5), 
            .O(readdata_c_15));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14883_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_552_i4_3_lut (.I0(n4568[203]), .I1(n4568[219]), .I2(address_c_0), 
            .I3(GND_net), .O(n4085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_552_i5_3_lut (.I0(n4568[204]), .I1(n4568[220]), .I2(address_c_0), 
            .I3(GND_net), .O(n4084));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_527_i15_4_lut (.I0(n4568[246]), .I1(\ootx_crc32_o[1] [14]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3690));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i15_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i19848_3_lut (.I0(n4551[3]), .I1(n4551[19]), .I2(address_c_0), 
            .I3(GND_net), .O(n24516));
    defparam i19848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14882_4_lut (.I0(n25864), .I1(n72), .I2(n3690), .I3(address_c_5), 
            .O(readdata_c_14));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14882_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i19849_3_lut (.I0(n4551[51]), .I1(n4551[67]), .I2(address_c_0), 
            .I3(GND_net), .O(n24517));
    defparam i19849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_527_i14_4_lut (.I0(n4568[245]), .I1(\ootx_crc32_o[1] [13]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3691));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i14_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i14881_4_lut (.I0(n25870), .I1(n72), .I2(n3691), .I3(address_c_5), 
            .O(readdata_c_13));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14881_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_527_i13_4_lut (.I0(n4568[244]), .I1(\ootx_crc32_o[1] [12]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3692));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i13_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i14880_4_lut (.I0(n25876), .I1(n72), .I2(n3692), .I3(address_c_5), 
            .O(readdata_c_12));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14880_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_527_i12_4_lut (.I0(n4568[243]), .I1(\ootx_crc32_o[1] [11]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3693));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i12_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i19867_3_lut (.I0(n4551[115]), .I1(n4551[123]), .I2(address_c_0), 
            .I3(GND_net), .O(n24535));
    defparam i19867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14879_4_lut (.I0(n25882), .I1(n72), .I2(n3693), .I3(address_c_5), 
            .O(readdata_c_11));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14879_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i19866_3_lut (.I0(n4551[83]), .I1(n4551[99]), .I2(address_c_0), 
            .I3(GND_net), .O(n24534));
    defparam i19866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19785_3_lut (.I0(n4551[2]), .I1(n4551[18]), .I2(address_c_0), 
            .I3(GND_net), .O(n24453));
    defparam i19785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19786_3_lut (.I0(n4551[50]), .I1(n4551[66]), .I2(address_c_0), 
            .I3(GND_net), .O(n24454));
    defparam i19786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19864_3_lut (.I0(n4551[114]), .I1(n4551[122]), .I2(address_c_0), 
            .I3(GND_net), .O(n24532));
    defparam i19864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19863_3_lut (.I0(n4551[82]), .I1(n4551[98]), .I2(address_c_0), 
            .I3(GND_net), .O(n24531));
    defparam i19863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_527_i11_4_lut (.I0(n4568[242]), .I1(\ootx_crc32_o[1] [10]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3694));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i11_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i14878_4_lut (.I0(n25888), .I1(n72), .I2(n3694), .I3(address_c_5), 
            .O(readdata_c_10));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14878_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_527_i10_4_lut (.I0(n4568[241]), .I1(\ootx_crc32_o[1] [9]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3695));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i10_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i14877_4_lut (.I0(n25204), .I1(n72), .I2(n3695), .I3(address_c_5), 
            .O(readdata_c_9));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14877_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 mux_527_i9_4_lut (.I0(n4568[240]), .I1(\ootx_crc32_o[1] [8]), 
            .I2(address_c_1), .I3(address_c_0), .O(n3696));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_527_i9_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i14876_4_lut (.I0(n25210), .I1(n72), .I2(n3696), .I3(address_c_5), 
            .O(readdata_c_8));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14876_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i14875_4_lut (.I0(n25216), .I1(n72), .I2(n25588), .I3(address_c_5), 
            .O(readdata_c_7));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14875_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14874_4_lut (.I0(n25228), .I1(n72), .I2(n25594), .I3(address_c_5), 
            .O(readdata_c_6));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14874_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14873_4_lut (.I0(n25240), .I1(n72), .I2(n25606), .I3(address_c_5), 
            .O(readdata_c_5));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14873_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14872_4_lut (.I0(n25246), .I1(n72), .I2(n25612), .I3(address_c_5), 
            .O(readdata_c_4));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14872_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i19788_3_lut (.I0(n4551[1]), .I1(n4551[17]), .I2(address_c_0), 
            .I3(GND_net), .O(n24456));
    defparam i19788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14871_4_lut (.I0(n25252), .I1(n72), .I2(n25624), .I3(address_c_5), 
            .O(readdata_c_3));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14871_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14870_4_lut (.I0(n25258), .I1(n72), .I2(n25630), .I3(address_c_5), 
            .O(readdata_c_2));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14870_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14869_4_lut (.I0(n25264), .I1(n72), .I2(n25636), .I3(address_c_5), 
            .O(readdata_c_1));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14869_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i14757_4_lut (.I0(n25564), .I1(n72), .I2(n25774), .I3(address_c_5), 
            .O(readdata_c_0));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14757_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i19789_3_lut (.I0(n4551[49]), .I1(n4551[65]), .I2(address_c_0), 
            .I3(GND_net), .O(n24457));
    defparam i19789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19861_3_lut (.I0(n4551[113]), .I1(n4551[121]), .I2(address_c_0), 
            .I3(GND_net), .O(n24529));
    defparam i19861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19860_3_lut (.I0(n4551[81]), .I1(n4551[97]), .I2(address_c_0), 
            .I3(GND_net), .O(n24528));
    defparam i19860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8000_3_lut_4_lut (.I0(n4551[172]), .I1(n1261), .I2(n22943), 
            .I3(n9513), .O(n12110));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8000_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7999_3_lut_4_lut (.I0(n4551[171]), .I1(n1262), .I2(n22943), 
            .I3(n9513), .O(n12109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7999_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19434_2_lut_3_lut (.I0(n13329), .I1(sensor_N_132), .I2(sensor_state), 
            .I3(GND_net), .O(n2));
    defparam i19434_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i7998_3_lut_4_lut (.I0(n4551[170]), .I1(n1263), .I2(n22943), 
            .I3(n9513), .O(n12108));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7998_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7997_3_lut_4_lut (.I0(n4551[169]), .I1(n1264), .I2(n22943), 
            .I3(n9513), .O(n12107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7997_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7996_3_lut_4_lut (.I0(n4551[168]), .I1(n1265), .I2(n22943), 
            .I3(n9513), .O(n12106));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7996_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19791_3_lut (.I0(sensor_signals_c_0), .I1(sensor_signals_c_1), 
            .I2(sensor_select[0]), .I3(GND_net), .O(n24459));
    defparam i19791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7995_3_lut_4_lut (.I0(n4551[167]), .I1(n1266), .I2(n22943), 
            .I3(n9513), .O(n12105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7995_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 sync_1__I_0_i1_2_lut (.I0(sync[0]), .I1(sync[1]), .I2(GND_net), 
            .I3(GND_net), .O(waitrequest_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(97[22:27])
    defparam sync_1__I_0_i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19792_3_lut (.I0(sensor_signals_c_2), .I1(sensor_signals_c_3), 
            .I2(sensor_select[0]), .I3(GND_net), .O(n24460));
    defparam i19792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7994_3_lut_4_lut (.I0(n4551[166]), .I1(n1267), .I2(n22943), 
            .I3(n9513), .O(n12104));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7994_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7993_3_lut_4_lut (.I0(n4551[165]), .I1(n1268), .I2(n22943), 
            .I3(n9513), .O(n12103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7993_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7992_3_lut_4_lut (.I0(n4551[164]), .I1(n1269), .I2(n22943), 
            .I3(n9513), .O(n12102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7992_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7991_3_lut_4_lut (.I0(n4551[163]), .I1(n1270), .I2(n22943), 
            .I3(n9513), .O(n12101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7991_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7990_3_lut_4_lut (.I0(n4551[162]), .I1(n1271), .I2(n22943), 
            .I3(n9513), .O(n12100));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7990_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19858_3_lut (.I0(sensor_signals_c_6), .I1(sensor_signals_c_7), 
            .I2(sensor_select[0]), .I3(GND_net), .O(n24526));
    defparam i19858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7989_3_lut_4_lut (.I0(n4551[161]), .I1(n1272), .I2(n22943), 
            .I3(n9513), .O(n12099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7989_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19857_3_lut (.I0(sensor_signals_c_4), .I1(sensor_signals_c_5), 
            .I2(sensor_select[0]), .I3(GND_net), .O(n24525));
    defparam i19857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7988_3_lut_4_lut (.I0(n4551[160]), .I1(n1273), .I2(n22943), 
            .I3(n9513), .O(n12098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7988_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7987_3_lut_4_lut (.I0(n4551[159]), .I1(n1274), .I2(n22943), 
            .I3(n9513), .O(n12097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7987_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7986_3_lut_4_lut (.I0(n4551[158]), .I1(n1275), .I2(n22943), 
            .I3(n9513), .O(n12096));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7986_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7985_3_lut_4_lut (.I0(n4551[157]), .I1(n1276), .I2(n22943), 
            .I3(n9513), .O(n12095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7985_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7984_3_lut_4_lut (.I0(n4551[156]), .I1(n1277), .I2(n22943), 
            .I3(n9513), .O(n12094));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7984_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7983_3_lut_4_lut (.I0(n4551[155]), .I1(n1278), .I2(n22943), 
            .I3(n9513), .O(n12093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7983_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7982_3_lut_4_lut (.I0(n4551[154]), .I1(n1279), .I2(n22943), 
            .I3(n9513), .O(n12092));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7982_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7981_3_lut_4_lut (.I0(n4551[153]), .I1(n1280), .I2(n22943), 
            .I3(n9513), .O(n12091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7981_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7980_3_lut_4_lut (.I0(n4551[152]), .I1(n1281), .I2(n22943), 
            .I3(n9513), .O(n12090));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7980_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7979_3_lut_4_lut (.I0(n4551[151]), .I1(n1282), .I2(n22943), 
            .I3(n9513), .O(n12089));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7979_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7978_3_lut_4_lut (.I0(n4551[150]), .I1(n1283), .I2(n22943), 
            .I3(n9513), .O(n12088));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7978_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19794_3_lut (.I0(n4551[256]), .I1(\ootx_crc32_o[0] [0]), .I2(address_c_0), 
            .I3(GND_net), .O(n24462));
    defparam i19794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7977_3_lut_4_lut (.I0(n4551[149]), .I1(n1284), .I2(n22943), 
            .I3(n9513), .O(n12087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7977_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19795_3_lut (.I0(n4568[0]), .I1(n4568[16]), .I2(address_c_0), 
            .I3(GND_net), .O(n24463));
    defparam i19795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7976_3_lut_4_lut (.I0(n4551[148]), .I1(n1285), .I2(n22943), 
            .I3(n9513), .O(n12086));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7976_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20406_4_lut (.I0(\ootx_crc32_o[0] [30]), .I1(n8917), .I2(n4568[46]), 
            .I3(address_c_1), .O(n24767));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20406_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7975_3_lut_4_lut (.I0(n4551[147]), .I1(n1286), .I2(n22943), 
            .I3(n9513), .O(n12085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7975_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7974_3_lut_4_lut (.I0(n4551[146]), .I1(n1287), .I2(n22943), 
            .I3(n9513), .O(n12084));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7974_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19855_3_lut (.I0(n4568[80]), .I1(n4568[96]), .I2(address_c_0), 
            .I3(GND_net), .O(n24523));
    defparam i19855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7973_3_lut_4_lut (.I0(n4551[145]), .I1(n1288), .I2(n22943), 
            .I3(n9513), .O(n12083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7973_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7972_3_lut_4_lut (.I0(n4551[144]), .I1(n1289), .I2(n22943), 
            .I3(n9513), .O(n12082));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7972_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_541_i31_4_lut (.I0(n4551[46]), .I1(n24767), .I2(address_c_4), 
            .I3(n13397), .O(n3912));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_541_i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i19854_3_lut (.I0(n4568[48]), .I1(n4568[64]), .I2(address_c_0), 
            .I3(GND_net), .O(n24522));
    defparam i19854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7971_3_lut_4_lut (.I0(n4551[143]), .I1(n1290), .I2(n22943), 
            .I3(n9513), .O(n12081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7971_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7970_3_lut_4_lut (.I0(n4551[142]), .I1(n1291), .I2(n22943), 
            .I3(n9513), .O(n12080));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7970_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19797_3_lut (.I0(n4551[0]), .I1(n4551[16]), .I2(address_c_0), 
            .I3(GND_net), .O(n24465));
    defparam i19797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14895_4_lut (.I0(n3912), .I1(n72), .I2(n24781), .I3(address_c_5), 
            .O(readdata_c_30));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i14895_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i7969_3_lut_4_lut (.I0(n4551[141]), .I1(n1292), .I2(n22943), 
            .I3(n9513), .O(n12079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7969_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7968_3_lut_4_lut (.I0(n4551[140]), .I1(n1293), .I2(n22943), 
            .I3(n9513), .O(n12078));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7968_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7967_3_lut_4_lut (.I0(n4551[139]), .I1(n1294), .I2(n22943), 
            .I3(n9513), .O(n12077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7967_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19798_3_lut (.I0(n4551[48]), .I1(n4551[64]), .I2(address_c_0), 
            .I3(GND_net), .O(n24466));
    defparam i19798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7966_3_lut_4_lut (.I0(n4551[138]), .I1(n1295), .I2(n22943), 
            .I3(n9513), .O(n12076));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7966_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7965_3_lut_4_lut (.I0(n4551[137]), .I1(n1296), .I2(n22943), 
            .I3(n9513), .O(n12075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7965_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19852_3_lut (.I0(n4551[112]), .I1(n4551[120]), .I2(address_c_0), 
            .I3(GND_net), .O(n24520));
    defparam i19852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7964_3_lut_4_lut (.I0(n4551[136]), .I1(n1297), .I2(n22943), 
            .I3(n9513), .O(n12074));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7964_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7963_3_lut_4_lut (.I0(n4551[135]), .I1(n1298), .I2(n22943), 
            .I3(n9513), .O(n12073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7963_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19851_3_lut (.I0(n4551[80]), .I1(n4551[96]), .I2(address_c_0), 
            .I3(GND_net), .O(n24519));
    defparam i19851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19800_3_lut (.I0(n4551[263]), .I1(\ootx_crc32_o[0] [7]), .I2(address_c_0), 
            .I3(GND_net), .O(n24468));
    defparam i19800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7962_3_lut_4_lut (.I0(n4551[134]), .I1(n1299), .I2(n22943), 
            .I3(n9513), .O(n12072));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7962_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7961_3_lut_4_lut (.I0(n4551[133]), .I1(n1300), .I2(n22943), 
            .I3(n9513), .O(n12071));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7961_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19801_3_lut (.I0(n4568[7]), .I1(n4568[23]), .I2(address_c_0), 
            .I3(GND_net), .O(n24469));
    defparam i19801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19750_3_lut (.I0(n4568[87]), .I1(n4568[103]), .I2(address_c_0), 
            .I3(GND_net), .O(n24418));
    defparam i19750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7960_3_lut_4_lut (.I0(n4551[132]), .I1(n1301), .I2(n22943), 
            .I3(n9513), .O(n12070));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7960_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7959_3_lut_4_lut (.I0(n4551[131]), .I1(n1302), .I2(n22943), 
            .I3(n9513), .O(n12069));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7959_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19749_3_lut (.I0(n4568[55]), .I1(n4568[71]), .I2(address_c_0), 
            .I3(GND_net), .O(n24417));
    defparam i19749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19818_3_lut (.I0(n4551[262]), .I1(\ootx_crc32_o[0] [6]), .I2(address_c_0), 
            .I3(GND_net), .O(n24486));
    defparam i19818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19819_3_lut (.I0(n4568[6]), .I1(n4568[22]), .I2(address_c_0), 
            .I3(GND_net), .O(n24487));
    defparam i19819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19726_3_lut (.I0(n4568[86]), .I1(n4568[102]), .I2(address_c_0), 
            .I3(GND_net), .O(n24394));
    defparam i19726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19725_3_lut (.I0(n4568[54]), .I1(n4568[70]), .I2(address_c_0), 
            .I3(GND_net), .O(n24393));
    defparam i19725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7958_3_lut_4_lut (.I0(n4551[130]), .I1(n1303), .I2(n22943), 
            .I3(n9513), .O(n12068));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7958_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7957_3_lut_4_lut (.I0(n4551[129]), .I1(n1304), .I2(n22943), 
            .I3(n9513), .O(n12067));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7957_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7956_3_lut_4_lut (.I0(n4551[128]), .I1(n1305), .I2(n22943), 
            .I3(n9513), .O(n12066));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7956_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7955_3_lut_4_lut (.I0(n4551[127]), .I1(n1306), .I2(n22943), 
            .I3(n9513), .O(n12065));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7955_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19821_3_lut (.I0(n4551[261]), .I1(\ootx_crc32_o[0] [5]), .I2(address_c_0), 
            .I3(GND_net), .O(n24489));
    defparam i19821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7954_3_lut_4_lut (.I0(n4551[126]), .I1(n1307), .I2(n22943), 
            .I3(n9513), .O(n12064));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7954_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19822_3_lut (.I0(n4568[5]), .I1(n4568[21]), .I2(address_c_0), 
            .I3(GND_net), .O(n24490));
    defparam i19822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7953_3_lut_4_lut (.I0(n4551[125]), .I1(n1308), .I2(n22943), 
            .I3(n9513), .O(n12063));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7953_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7952_3_lut_4_lut (.I0(n4551[124]), .I1(n1309), .I2(n22943), 
            .I3(n9513), .O(n12062));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7952_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7951_3_lut_4_lut (.I0(n4551[123]), .I1(n1310), .I2(n22943), 
            .I3(n9513), .O(n12061));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7951_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7950_3_lut_4_lut (.I0(n4551[122]), .I1(n1311), .I2(n22943), 
            .I3(n9513), .O(n12060));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7950_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7949_3_lut_4_lut (.I0(n4551[121]), .I1(n1312), .I2(n22943), 
            .I3(n9513), .O(n12059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7949_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7948_3_lut_4_lut (.I0(n4551[120]), .I1(n1313), .I2(n22943), 
            .I3(n9513), .O(n12058));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7948_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19699_3_lut (.I0(n4568[85]), .I1(n4568[101]), .I2(address_c_0), 
            .I3(GND_net), .O(n24367));
    defparam i19699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14733_2_lut_3_lut (.I0(n2679), .I1(n9200), .I2(ootx_payloads_N_1699[30]), 
            .I3(GND_net), .O(ootx_payloads_N_1698));
    defparam i14733_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i7947_3_lut_4_lut (.I0(n4551[119]), .I1(n1314), .I2(n22943), 
            .I3(n9513), .O(n12057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7947_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19698_3_lut (.I0(n4568[53]), .I1(n4568[69]), .I2(address_c_0), 
            .I3(GND_net), .O(n24366));
    defparam i19698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7946_3_lut_4_lut (.I0(n4551[118]), .I1(n1315), .I2(n22943), 
            .I3(n9513), .O(n12056));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7946_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7945_3_lut_4_lut (.I0(n4551[117]), .I1(n1316), .I2(n22943), 
            .I3(n9513), .O(n12055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7945_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7944_3_lut_4_lut (.I0(n4551[116]), .I1(n1317), .I2(n22943), 
            .I3(n9513), .O(n12054));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7944_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7943_3_lut_4_lut (.I0(n4551[115]), .I1(n1318), .I2(n22943), 
            .I3(n9513), .O(n12053));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7943_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7942_3_lut_4_lut (.I0(n4551[114]), .I1(n1319), .I2(n22943), 
            .I3(n9513), .O(n12052));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7942_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7941_3_lut_4_lut (.I0(n4551[113]), .I1(n1320), .I2(n22943), 
            .I3(n9513), .O(n12051));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7941_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7940_3_lut_4_lut (.I0(n4551[112]), .I1(n1321), .I2(n22943), 
            .I3(n9513), .O(n12050));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7940_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19824_3_lut (.I0(n4551[260]), .I1(\ootx_crc32_o[0] [4]), .I2(address_c_0), 
            .I3(GND_net), .O(n24492));
    defparam i19824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7939_3_lut_4_lut (.I0(n4551[111]), .I1(n1322), .I2(n22943), 
            .I3(n9513), .O(n12049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7939_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19825_3_lut (.I0(n4568[4]), .I1(n4568[20]), .I2(address_c_0), 
            .I3(GND_net), .O(n24493));
    defparam i19825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7938_3_lut_4_lut (.I0(n4551[110]), .I1(n1323), .I2(n22943), 
            .I3(n9513), .O(n12048));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7938_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19696_3_lut (.I0(n4568[84]), .I1(n4568[100]), .I2(address_c_0), 
            .I3(GND_net), .O(n24364));
    defparam i19696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7937_3_lut_4_lut (.I0(n4551[109]), .I1(n1324), .I2(n22943), 
            .I3(n9513), .O(n12047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7937_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19695_3_lut (.I0(n4568[52]), .I1(n4568[68]), .I2(address_c_0), 
            .I3(GND_net), .O(n24363));
    defparam i19695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7936_3_lut_4_lut (.I0(n4551[108]), .I1(n1325), .I2(n22943), 
            .I3(n9513), .O(n12046));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7936_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7935_3_lut_4_lut (.I0(n4551[107]), .I1(n1326), .I2(n22943), 
            .I3(n9513), .O(n12045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7935_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7934_3_lut_4_lut (.I0(n4551[106]), .I1(n1327), .I2(n22943), 
            .I3(n9513), .O(n12044));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7934_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7933_3_lut_4_lut (.I0(n4551[105]), .I1(n1328), .I2(n22943), 
            .I3(n9513), .O(n12043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7933_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19827_3_lut (.I0(n4551[259]), .I1(\ootx_crc32_o[0] [3]), .I2(address_c_0), 
            .I3(GND_net), .O(n24495));
    defparam i19827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7932_3_lut_4_lut (.I0(n4551[104]), .I1(n1329), .I2(n22943), 
            .I3(n9513), .O(n12042));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7932_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7931_3_lut_4_lut (.I0(n4551[103]), .I1(n1330), .I2(n22943), 
            .I3(n9513), .O(n12041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7931_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7930_3_lut_4_lut (.I0(n4551[102]), .I1(n1331), .I2(n22943), 
            .I3(n9513), .O(n12040));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7930_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19828_3_lut (.I0(n4568[3]), .I1(n4568[19]), .I2(address_c_0), 
            .I3(GND_net), .O(n24496));
    defparam i19828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7929_3_lut_4_lut (.I0(n4551[101]), .I1(n1332), .I2(n22943), 
            .I3(n9513), .O(n12039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7929_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7928_3_lut_4_lut (.I0(n4551[100]), .I1(n1333), .I2(n22943), 
            .I3(n9513), .O(n12038));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7928_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7927_3_lut_4_lut (.I0(n4551[99]), .I1(n1334), .I2(n22943), 
            .I3(n9513), .O(n12037));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7927_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7926_3_lut_4_lut (.I0(n4551[98]), .I1(n1335), .I2(n22943), 
            .I3(n9513), .O(n12036));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7926_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7925_3_lut_4_lut (.I0(n4551[97]), .I1(n1336), .I2(n22943), 
            .I3(n9513), .O(n12035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7925_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19648_3_lut (.I0(n4568[83]), .I1(n4568[99]), .I2(address_c_0), 
            .I3(GND_net), .O(n24316));
    defparam i19648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7924_3_lut_4_lut (.I0(n4551[96]), .I1(n1337), .I2(n22943), 
            .I3(n9513), .O(n12034));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7924_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7923_3_lut_4_lut (.I0(n4551[95]), .I1(n1338), .I2(n22943), 
            .I3(n9513), .O(n12033));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7923_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7922_3_lut_4_lut (.I0(n4551[94]), .I1(n1339), .I2(n22943), 
            .I3(n9513), .O(n12032));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7922_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7921_3_lut_4_lut (.I0(n4551[93]), .I1(n1340), .I2(n22943), 
            .I3(n9513), .O(n12031));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7921_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7920_3_lut_4_lut (.I0(n4551[92]), .I1(n1341), .I2(n22943), 
            .I3(n9513), .O(n12030));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7920_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19647_3_lut (.I0(n4568[51]), .I1(n4568[67]), .I2(address_c_0), 
            .I3(GND_net), .O(n24315));
    defparam i19647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7919_3_lut_4_lut (.I0(n4551[91]), .I1(n1342), .I2(n22943), 
            .I3(n9513), .O(n12029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7919_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19830_3_lut (.I0(n4551[258]), .I1(\ootx_crc32_o[0] [2]), .I2(address_c_0), 
            .I3(GND_net), .O(n24498));
    defparam i19830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7918_3_lut_4_lut (.I0(n4551[90]), .I1(n1343), .I2(n22943), 
            .I3(n9513), .O(n12028));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7918_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19831_3_lut (.I0(n4568[2]), .I1(n4568[18]), .I2(address_c_0), 
            .I3(GND_net), .O(n24499));
    defparam i19831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7917_3_lut_4_lut (.I0(n4551[89]), .I1(n1344), .I2(n22943), 
            .I3(n9513), .O(n12027));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7917_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7916_3_lut_4_lut (.I0(n4551[88]), .I1(n1345), .I2(n22943), 
            .I3(n9513), .O(n12026));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7916_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7915_3_lut_4_lut (.I0(n4551[87]), .I1(n1346), .I2(n22943), 
            .I3(n9513), .O(n12025));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7915_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(n9200), .I1(ootx_payloads_N_1699[30]), 
            .I2(GND_net), .I3(GND_net), .O(n2680));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'heeee;
    SB_LUT4 i7914_3_lut_4_lut (.I0(n4551[86]), .I1(n1347), .I2(n22943), 
            .I3(n9513), .O(n12024));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7914_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7913_3_lut_4_lut (.I0(n4551[85]), .I1(n1348), .I2(n22943), 
            .I3(n9513), .O(n12023));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7913_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7912_3_lut_4_lut (.I0(n4551[84]), .I1(n1349), .I2(n22943), 
            .I3(n9513), .O(n12022));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7912_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7911_3_lut_4_lut (.I0(n4551[83]), .I1(n1350), .I2(n22943), 
            .I3(n9513), .O(n12021));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7911_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7910_3_lut_4_lut (.I0(n4551[82]), .I1(n1351), .I2(n22943), 
            .I3(n9513), .O(n12020));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7910_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7909_3_lut_4_lut (.I0(n4551[81]), .I1(n1352), .I2(n22943), 
            .I3(n9513), .O(n12019));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7909_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7908_3_lut_4_lut (.I0(n4551[80]), .I1(n1353), .I2(n22943), 
            .I3(n9513), .O(n12018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7908_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7907_3_lut_4_lut (.I0(n4551[79]), .I1(n1354), .I2(n22943), 
            .I3(n9513), .O(n12017));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7907_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7906_3_lut_4_lut (.I0(n4551[78]), .I1(n1355), .I2(n22943), 
            .I3(n9513), .O(n12016));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7906_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19645_3_lut (.I0(n4568[82]), .I1(n4568[98]), .I2(address_c_0), 
            .I3(GND_net), .O(n24313));
    defparam i19645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19644_3_lut (.I0(n4568[50]), .I1(n4568[66]), .I2(address_c_0), 
            .I3(GND_net), .O(n24312));
    defparam i19644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_425_i10_4_lut (.I0(ootx_payloads_N_1730[0]), .I1(ootx_payloads_N_1730[1]), 
            .I2(ootx_payloads_N_1699[4]), .I3(ootx_payloads_N_1699[3]), 
            .O(n10));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i10_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i7905_3_lut_4_lut (.I0(n4551[77]), .I1(n1356), .I2(n22943), 
            .I3(n9513), .O(n12015));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7905_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7904_3_lut_4_lut (.I0(n4551[76]), .I1(n1357), .I2(n22943), 
            .I3(n9513), .O(n12014));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7904_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1044 (.I0(ootx_payloads_N_1744[0]), .I1(n2679), 
            .I2(n9200), .I3(ootx_payloads_N_1699[30]), .O(n30_adj_2286));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1044.LUT_INIT = 16'haaae;
    SB_LUT4 i19833_3_lut (.I0(n4551[257]), .I1(\ootx_crc32_o[0] [1]), .I2(address_c_0), 
            .I3(GND_net), .O(n24501));
    defparam i19833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7903_3_lut_4_lut (.I0(n4551[75]), .I1(n1358), .I2(n22943), 
            .I3(n9513), .O(n12013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7903_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7902_3_lut_4_lut (.I0(n4551[74]), .I1(n1359), .I2(n22943), 
            .I3(n9513), .O(n12012));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7902_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7901_3_lut_4_lut (.I0(n4551[73]), .I1(n1360), .I2(n22943), 
            .I3(n9513), .O(n12011));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7901_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7900_3_lut_4_lut (.I0(n4551[72]), .I1(n1361), .I2(n22943), 
            .I3(n9513), .O(n12010));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7900_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7899_3_lut_4_lut (.I0(n4551[71]), .I1(n1362), .I2(n22943), 
            .I3(n9513), .O(n12009));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7899_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7898_3_lut_4_lut (.I0(n4551[70]), .I1(n1363), .I2(n22943), 
            .I3(n9513), .O(n12008));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7898_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i12_3_lut (.I0(n10), .I1(ootx_payloads_N_1730[2]), 
            .I2(ootx_payloads_N_1699[5]), .I3(GND_net), .O(n12));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i19834_3_lut (.I0(n4568[1]), .I1(n4568[17]), .I2(address_c_0), 
            .I3(GND_net), .O(n24502));
    defparam i19834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7897_3_lut_4_lut (.I0(n4551[69]), .I1(n1364), .I2(n22943), 
            .I3(n9513), .O(n12007));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7897_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7896_3_lut_4_lut (.I0(n4551[68]), .I1(n1365), .I2(n22943), 
            .I3(n9513), .O(n12006));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7896_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7895_3_lut_4_lut (.I0(n4551[67]), .I1(n1366), .I2(n22943), 
            .I3(n9513), .O(n12005));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7895_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19642_3_lut (.I0(n4568[81]), .I1(n4568[97]), .I2(address_c_0), 
            .I3(GND_net), .O(n24310));
    defparam i19642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20416_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[179]), .O(n24831));
    defparam i20416_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i20415_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[181]), .O(n24801));
    defparam i20415_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i7894_3_lut_4_lut (.I0(n4551[66]), .I1(n1367), .I2(n22943), 
            .I3(n9513), .O(n12004));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7894_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7893_3_lut_4_lut (.I0(n4551[65]), .I1(n1368), .I2(n22943), 
            .I3(n9513), .O(n12003));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7893_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19641_3_lut (.I0(n4568[49]), .I1(n4568[65]), .I2(address_c_0), 
            .I3(GND_net), .O(n24309));
    defparam i19641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19836_3_lut (.I0(n4551[7]), .I1(n4551[23]), .I2(address_c_0), 
            .I3(GND_net), .O(n24504));
    defparam i19836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7892_3_lut_4_lut (.I0(n4551[64]), .I1(n1369), .I2(n22943), 
            .I3(n9513), .O(n12002));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7892_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7891_3_lut_4_lut (.I0(n4551[63]), .I1(n1370), .I2(n22943), 
            .I3(n9513), .O(n12001));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7891_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7890_3_lut_4_lut (.I0(n4551[62]), .I1(n1371), .I2(n22943), 
            .I3(n9513), .O(n12000));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7890_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19837_3_lut (.I0(n4551[55]), .I1(n4551[71]), .I2(address_c_0), 
            .I3(GND_net), .O(n24505));
    defparam i19837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7889_3_lut_4_lut (.I0(n4551[61]), .I1(n1372), .I2(n22943), 
            .I3(n9513), .O(n11999));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7889_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7888_3_lut_4_lut (.I0(n4551[60]), .I1(n1373), .I2(n22943), 
            .I3(n9513), .O(n11998));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7888_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7887_3_lut_4_lut (.I0(n4551[59]), .I1(n1374), .I2(n22943), 
            .I3(n9513), .O(n11997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7887_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7886_3_lut_4_lut (.I0(n4551[58]), .I1(n1375), .I2(n22943), 
            .I3(n9513), .O(n11996));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7886_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7885_3_lut_4_lut (.I0(n4551[57]), .I1(n1376), .I2(n22943), 
            .I3(n9513), .O(n11995));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7885_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7884_3_lut_4_lut (.I0(n4551[56]), .I1(n1377), .I2(n22943), 
            .I3(n9513), .O(n11994));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7884_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7883_3_lut_4_lut (.I0(n4551[55]), .I1(n1378), .I2(n22943), 
            .I3(n9513), .O(n11993));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7883_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i14_3_lut (.I0(n12), .I1(ootx_payloads_N_1730[3]), 
            .I2(ootx_payloads_N_1699[6]), .I3(GND_net), .O(n14));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7882_3_lut_4_lut (.I0(n4551[54]), .I1(n1379), .I2(n22943), 
            .I3(n9513), .O(n11992));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7882_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7881_3_lut_4_lut (.I0(n4551[53]), .I1(n1380), .I2(n22943), 
            .I3(n9513), .O(n11991));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7881_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7880_3_lut_4_lut (.I0(n4551[52]), .I1(n1381), .I2(n22943), 
            .I3(n9513), .O(n11990));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7880_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19639_3_lut (.I0(n4551[119]), .I1(n4551[127]), .I2(address_c_0), 
            .I3(GND_net), .O(n24307));
    defparam i19639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_425_i16_3_lut (.I0(n14), .I1(ootx_payloads_N_1730[4]), 
            .I2(ootx_payloads_N_1699[7]), .I3(GND_net), .O(n16));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i20452_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[182]), .O(n24826));
    defparam i20452_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 LessThan_425_i18_3_lut (.I0(n16), .I1(ootx_payloads_N_1730[5]), 
            .I2(ootx_payloads_N_1699[8]), .I3(GND_net), .O(n18));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7879_3_lut_4_lut (.I0(n4551[51]), .I1(n1382), .I2(n22943), 
            .I3(n9513), .O(n11989));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7879_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7878_3_lut_4_lut (.I0(n4551[50]), .I1(n1383), .I2(n22943), 
            .I3(n9513), .O(n11988));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7878_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7877_3_lut_4_lut (.I0(n4551[49]), .I1(n1384), .I2(n22943), 
            .I3(n9513), .O(n11987));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7877_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19638_3_lut (.I0(n4551[87]), .I1(n4551[103]), .I2(address_c_0), 
            .I3(GND_net), .O(n24306));
    defparam i19638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_425_i20_3_lut (.I0(n18), .I1(ootx_payloads_N_1730[6]), 
            .I2(ootx_payloads_N_1699[9]), .I3(GND_net), .O(n20));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7876_3_lut_4_lut (.I0(n4551[48]), .I1(n1385), .I2(n22943), 
            .I3(n9513), .O(n11986));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7876_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_552_i6_3_lut (.I0(n4568[205]), .I1(n4568[221]), .I2(address_c_0), 
            .I3(GND_net), .O(n4083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7875_3_lut_4_lut (.I0(n4551[47]), .I1(n1386), .I2(n22943), 
            .I3(n9513), .O(n11985));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7875_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7874_3_lut_4_lut (.I0(n4551[46]), .I1(n1387), .I2(n22943), 
            .I3(n9513), .O(n11984));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7874_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i22_3_lut (.I0(n20), .I1(ootx_payloads_N_1730[7]), 
            .I2(ootx_payloads_N_1699[10]), .I3(GND_net), .O(n22));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7873_3_lut_4_lut (.I0(n4551[45]), .I1(n1388), .I2(n22943), 
            .I3(n9513), .O(n11983));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7873_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7872_3_lut_4_lut (.I0(n4551[44]), .I1(n1389), .I2(n22943), 
            .I3(n9513), .O(n11982));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7872_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20417_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[178]), .O(n24833));
    defparam i20417_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i19839_3_lut (.I0(n4551[6]), .I1(n4551[22]), .I2(address_c_0), 
            .I3(GND_net), .O(n24507));
    defparam i19839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20414_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[183]), .O(n24799));
    defparam i20414_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 LessThan_425_i24_3_lut (.I0(n22), .I1(ootx_payloads_N_1730[8]), 
            .I2(ootx_payloads_N_1699[11]), .I3(GND_net), .O(n24));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i20284_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[177]), .O(n24797));
    defparam i20284_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i20454_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[180]), .O(n24795));
    defparam i20454_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i20418_2_lut_3_lut_4_lut (.I0(n4702), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4568[176]), .O(n24617));
    defparam i20418_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i7871_3_lut_4_lut (.I0(n4551[43]), .I1(n1390), .I2(n22943), 
            .I3(n9513), .O(n11981));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7871_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7870_3_lut_4_lut (.I0(n4551[42]), .I1(n1391), .I2(n22943), 
            .I3(n9513), .O(n11980));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7870_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7869_3_lut_4_lut (.I0(n4551[41]), .I1(n1392), .I2(n22943), 
            .I3(n9513), .O(n11979));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7869_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7868_3_lut_4_lut (.I0(n4551[40]), .I1(n1393), .I2(n22943), 
            .I3(n9513), .O(n11978));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7868_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7867_3_lut_4_lut (.I0(n4551[39]), .I1(n1394), .I2(n22943), 
            .I3(n9513), .O(n11977));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7867_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19840_3_lut (.I0(n4551[54]), .I1(n4551[70]), .I2(address_c_0), 
            .I3(GND_net), .O(n24508));
    defparam i19840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7866_3_lut_4_lut (.I0(n4551[38]), .I1(n1395), .I2(n22943), 
            .I3(n9513), .O(n11976));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7866_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19615_3_lut (.I0(n4551[118]), .I1(n4551[126]), .I2(address_c_0), 
            .I3(GND_net), .O(n24283));
    defparam i19615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7865_3_lut_4_lut (.I0(n4551[37]), .I1(n1396), .I2(n22943), 
            .I3(n9513), .O(n11975));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7865_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19614_3_lut (.I0(n4551[86]), .I1(n4551[102]), .I2(address_c_0), 
            .I3(GND_net), .O(n24282));
    defparam i19614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7864_3_lut_4_lut (.I0(n4551[36]), .I1(n1397), .I2(n22943), 
            .I3(n9513), .O(n11974));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7864_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7863_3_lut_4_lut (.I0(n4551[35]), .I1(n1398), .I2(n22943), 
            .I3(n9513), .O(n11973));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7863_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7862_3_lut_4_lut (.I0(n4551[34]), .I1(n1399), .I2(n22943), 
            .I3(n9513), .O(n11972));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7862_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i26_3_lut (.I0(n24), .I1(ootx_payloads_N_1730[9]), 
            .I2(ootx_payloads_N_1699[12]), .I3(GND_net), .O(n26));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7861_3_lut_4_lut (.I0(n4551[33]), .I1(n1400), .I2(n22943), 
            .I3(n9513), .O(n11971));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7861_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i28_3_lut (.I0(n26), .I1(ootx_payloads_N_1730[10]), 
            .I2(ootx_payloads_N_1699[13]), .I3(GND_net), .O(n28));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7860_3_lut_4_lut (.I0(n4551[32]), .I1(n1401), .I2(n22943), 
            .I3(n9513), .O(n11970));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7860_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i30_3_lut (.I0(n28), .I1(ootx_payloads_N_1730[11]), 
            .I2(ootx_payloads_N_1699[14]), .I3(GND_net), .O(n30));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7859_3_lut_4_lut (.I0(n4551[31]), .I1(n1402), .I2(n22943), 
            .I3(n9513), .O(n11969));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7859_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7858_3_lut_4_lut (.I0(n4551[30]), .I1(n1403), .I2(n22943), 
            .I3(n9513), .O(n11968));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7858_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 LessThan_425_i32_3_lut (.I0(n30), .I1(ootx_payloads_N_1730[12]), 
            .I2(ootx_payloads_N_1699[15]), .I3(GND_net), .O(n2679));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[10:80])
    defparam LessThan_425_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7857_3_lut_4_lut (.I0(n4551[29]), .I1(n1404), .I2(n22943), 
            .I3(n9513), .O(n11967));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7857_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7856_3_lut_4_lut (.I0(n4551[28]), .I1(n1405), .I2(n22943), 
            .I3(n9513), .O(n11966));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7856_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7855_3_lut_4_lut (.I0(n4551[27]), .I1(n1406), .I2(n22943), 
            .I3(n9513), .O(n11965));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7855_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7854_3_lut_4_lut (.I0(n4551[26]), .I1(n1407), .I2(n22943), 
            .I3(n9513), .O(n11964));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7854_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7853_3_lut_4_lut (.I0(n4551[25]), .I1(n1408), .I2(n22943), 
            .I3(n9513), .O(n11963));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7853_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7852_3_lut_4_lut (.I0(n4551[24]), .I1(n1409), .I2(n22943), 
            .I3(n9513), .O(n11962));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7852_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7851_3_lut_4_lut (.I0(n4551[23]), .I1(n1410), .I2(n22943), 
            .I3(n9513), .O(n11961));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7851_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19845_3_lut (.I0(n4551[4]), .I1(n4551[20]), .I2(address_c_0), 
            .I3(GND_net), .O(n24513));
    defparam i19845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19846_3_lut (.I0(n4551[52]), .I1(n4551[68]), .I2(address_c_0), 
            .I3(GND_net), .O(n24514));
    defparam i19846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7850_3_lut_4_lut (.I0(n4551[22]), .I1(n1411), .I2(n22943), 
            .I3(n9513), .O(n11960));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7850_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7849_3_lut_4_lut (.I0(n4551[21]), .I1(n1412), .I2(n22943), 
            .I3(n9513), .O(n11959));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7849_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i19480_3_lut (.I0(n4551[116]), .I1(n4551[124]), .I2(address_c_0), 
            .I3(GND_net), .O(n24148));
    defparam i19480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19479_3_lut (.I0(n4551[84]), .I1(n4551[100]), .I2(address_c_0), 
            .I3(GND_net), .O(n24147));
    defparam i19479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_552_i7_3_lut (.I0(n4568[206]), .I1(n4568[222]), .I2(address_c_0), 
            .I3(GND_net), .O(n4082));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_553_i2_3_lut (.I0(n4551[129]), .I1(n4551[145]), .I2(address_c_0), 
            .I3(GND_net), .O(n4104));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7848_3_lut_4_lut (.I0(n4551[20]), .I1(n1413), .I2(n22943), 
            .I3(n9513), .O(n11958));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7848_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7847_3_lut_4_lut (.I0(n4551[19]), .I1(n1414), .I2(n22943), 
            .I3(n9513), .O(n11957));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7847_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20282_4_lut (.I0(\ootx_crc32_o[0] [20]), .I1(n7584), .I2(n4568[36]), 
            .I3(address_c_1), .O(n24731));
    defparam i20282_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7846_3_lut_4_lut (.I0(n4551[18]), .I1(n1415), .I2(n22943), 
            .I3(n9513), .O(n11956));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7846_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7845_3_lut_4_lut (.I0(n4551[17]), .I1(n1416), .I2(n22943), 
            .I3(n9513), .O(n11955));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7845_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7844_3_lut_4_lut (.I0(n4551[16]), .I1(n1417), .I2(n22943), 
            .I3(n9513), .O(n11954));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7844_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7843_3_lut_4_lut (.I0(n4551[15]), .I1(n1418), .I2(n22943), 
            .I3(n9513), .O(n11953));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7843_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_553_i5_3_lut (.I0(n4551[132]), .I1(n4551[148]), .I2(address_c_0), 
            .I3(GND_net), .O(n4101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20423_4_lut (.I0(\ootx_crc32_o[0] [17]), .I1(n7584), .I2(n4568[33]), 
            .I3(address_c_1), .O(n24729));
    defparam i20423_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7842_3_lut_4_lut (.I0(n4551[14]), .I1(n1419), .I2(n22943), 
            .I3(n9513), .O(n11952));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7842_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7841_3_lut_4_lut (.I0(n4551[13]), .I1(n1420), .I2(n22943), 
            .I3(n9513), .O(n11951));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7841_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_553_i6_3_lut (.I0(n4551[133]), .I1(n4551[149]), .I2(address_c_0), 
            .I3(GND_net), .O(n4100));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_553_i7_3_lut (.I0(n4551[134]), .I1(n4551[150]), .I2(address_c_0), 
            .I3(GND_net), .O(n4099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7840_3_lut_4_lut (.I0(n4551[12]), .I1(n1421), .I2(n22943), 
            .I3(n9513), .O(n11950));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7840_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7839_3_lut_4_lut (.I0(n4551[11]), .I1(n1422), .I2(n22943), 
            .I3(n9513), .O(n11949));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7839_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7838_3_lut_4_lut (.I0(n4551[10]), .I1(n1423), .I2(n22943), 
            .I3(n9513), .O(n11948));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7838_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7837_3_lut_4_lut (.I0(n4551[9]), .I1(n1424), .I2(n22943), 
            .I3(n9513), .O(n11947));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7837_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7836_3_lut_4_lut (.I0(n4551[8]), .I1(n1425), .I2(n22943), 
            .I3(n9513), .O(n11946));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7836_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7835_3_lut_4_lut (.I0(n4551[7]), .I1(n1426), .I2(n22943), 
            .I3(n9513), .O(n11945));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7835_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7834_3_lut_4_lut (.I0(n4551[6]), .I1(n1427), .I2(n22943), 
            .I3(n9513), .O(n11944));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7834_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7833_3_lut_4_lut (.I0(n4551[5]), .I1(n1428), .I2(n22943), 
            .I3(n9513), .O(n11943));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7833_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7832_3_lut_4_lut (.I0(n4551[4]), .I1(n1429), .I2(n22943), 
            .I3(n9513), .O(n11942));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7832_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7831_3_lut_4_lut (.I0(n4551[3]), .I1(n1430), .I2(n22943), 
            .I3(n9513), .O(n11941));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7831_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7830_3_lut_4_lut (.I0(n4551[2]), .I1(n1431), .I2(n22943), 
            .I3(n9513), .O(n11940));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7830_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i7829_3_lut_4_lut (.I0(n4551[1]), .I1(n1432), .I2(n22943), 
            .I3(n9513), .O(n11939));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i7829_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20285_4_lut (.I0(\ootx_crc32_o[0] [23]), .I1(n7584), .I2(n4568[39]), 
            .I3(address_c_1), .O(n24798));
    defparam i20285_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20331_2_lut_3_lut (.I0(sensor_state), .I1(n13329), .I2(sensor_N_132), 
            .I3(GND_net), .O(n24692));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    defparam i20331_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20428_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [29]), 
            .I3(GND_net), .O(n24780));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20428_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20439_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [28]), 
            .I3(GND_net), .O(n24779));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20439_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20430_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [27]), 
            .I3(GND_net), .O(n24777));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20430_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20431_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [26]), 
            .I3(GND_net), .O(n24776));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20431_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20432_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [25]), 
            .I3(GND_net), .O(n24775));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20432_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20398_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [24]), 
            .I3(GND_net), .O(n24774));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20398_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6906_3_lut_4_lut (.I0(n4551[0]), .I1(n1433), .I2(n22943), 
            .I3(n9513), .O(n11016));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i6906_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20434_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [23]), 
            .I3(GND_net), .O(n24772));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20434_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20270_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [22]), 
            .I3(GND_net), .O(n24639));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20270_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20435_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [21]), 
            .I3(GND_net), .O(n24771));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20435_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20277_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [20]), 
            .I3(GND_net), .O(n24642));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20277_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20446_4_lut (.I0(\ootx_crc32_o[0] [21]), .I1(n7584), .I2(n4568[37]), 
            .I3(address_c_1), .O(n24800));
    defparam i20446_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i8_3_lut (.I0(n4568[207]), .I1(n4568[223]), .I2(address_c_0), 
            .I3(GND_net), .O(n4081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20436_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [19]), 
            .I3(GND_net), .O(n24770));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20436_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20366_4_lut (.I0(n4568[136]), .I1(address_c_1), .I2(n4568[152]), 
            .I3(address_c_0), .O(n24628));
    defparam i20366_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut (.I0(address_c_3), .I1(address_c_2), .I2(address_c_0), 
            .I3(GND_net), .O(n50_adj_2283));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i20437_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [18]), 
            .I3(GND_net), .O(n24769));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20437_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20276_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [17]), 
            .I3(GND_net), .O(n24643));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20276_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_552_i9_3_lut (.I0(n4568[208]), .I1(n4568[224]), .I2(address_c_0), 
            .I3(GND_net), .O(n4080));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20408_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [31]), 
            .I3(GND_net), .O(n24783));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20408_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20407_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [16]), 
            .I3(GND_net), .O(n24768));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20407_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20427_2_lut_3_lut (.I0(address_c_0), .I1(address_c_1), .I2(\ootx_crc32_o[1] [30]), 
            .I3(GND_net), .O(n24781));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam i20427_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20421_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[179]), .O(n24656));
    defparam i20421_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_adj_1045 (.I0(address_c_2), .I1(address_c_3), 
            .I2(address_c_0), .I3(GND_net), .O(n8917));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i1_2_lut_3_lut_adj_1045.LUT_INIT = 16'h1010;
    SB_LUT4 i20450_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[182]), .O(n24825));
    defparam i20450_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i20420_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[181]), .O(n24725));
    defparam i20420_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_3_lut_4_lut (.I0(address_c_2), .I1(address_c_3), .I2(address_c_5), 
            .I3(address_c_4), .O(n72));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(43[14:21])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf0e0;
    SB_LUT4 i20422_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[178]), .O(n24654));
    defparam i20422_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i20419_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[183]), .O(n24727));
    defparam i20419_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i20458_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[177]), .O(n24796));
    defparam i20458_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i20382_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[180]), .O(n24794));
    defparam i20382_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i20424_2_lut_3_lut_4_lut (.I0(n4673), .I1(address_c_1), .I2(address_c_2), 
            .I3(n4551[176]), .O(n24635));
    defparam i20424_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i8091_3_lut_4_lut (.I0(n4551[263]), .I1(n1170), .I2(n22943), 
            .I3(n9513), .O(n12201));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8091_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8090_3_lut_4_lut (.I0(n4551[262]), .I1(n1171), .I2(n22943), 
            .I3(n9513), .O(n12200));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8090_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20367_4_lut (.I0(n4568[137]), .I1(address_c_1), .I2(n4568[153]), 
            .I3(address_c_0), .O(n24627));
    defparam i20367_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_552_i10_3_lut (.I0(n4568[209]), .I1(n4568[225]), .I2(address_c_0), 
            .I3(GND_net), .O(n4079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_552_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8089_3_lut_4_lut (.I0(n4551[261]), .I1(n1172), .I2(n22943), 
            .I3(n9513), .O(n12199));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8089_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8088_3_lut_4_lut (.I0(n4551[260]), .I1(n1173), .I2(n22943), 
            .I3(n9513), .O(n12198));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8088_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8087_3_lut_4_lut (.I0(n4551[259]), .I1(n1174), .I2(n22943), 
            .I3(n9513), .O(n12197));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8087_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8086_3_lut_4_lut (.I0(n4551[258]), .I1(n1175), .I2(n22943), 
            .I3(n9513), .O(n12196));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8086_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8085_3_lut_4_lut (.I0(n4551[257]), .I1(n1176), .I2(n22943), 
            .I3(n9513), .O(n12195));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8085_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8084_3_lut_4_lut (.I0(n4551[256]), .I1(n1177), .I2(n22943), 
            .I3(n9513), .O(n12194));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8084_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8083_3_lut_4_lut (.I0(n4551[255]), .I1(n1178), .I2(n22943), 
            .I3(n9513), .O(n12193));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8083_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8082_3_lut_4_lut (.I0(n4551[254]), .I1(n1179), .I2(n22943), 
            .I3(n9513), .O(n12192));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8082_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8081_3_lut_4_lut (.I0(n4551[253]), .I1(n1180), .I2(n22943), 
            .I3(n9513), .O(n12191));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8081_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8080_3_lut_4_lut (.I0(n4551[252]), .I1(n1181), .I2(n22943), 
            .I3(n9513), .O(n12190));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8080_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8079_3_lut_4_lut (.I0(n4551[251]), .I1(n1182), .I2(n22943), 
            .I3(n9513), .O(n12189));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8079_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8078_3_lut_4_lut (.I0(n4551[250]), .I1(n1183), .I2(n22943), 
            .I3(n9513), .O(n12188));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8078_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8077_3_lut_4_lut (.I0(n4551[249]), .I1(n1184), .I2(n22943), 
            .I3(n9513), .O(n12187));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8077_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8076_3_lut_4_lut (.I0(n4551[248]), .I1(n1185), .I2(n22943), 
            .I3(n9513), .O(n12186));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8076_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8075_3_lut_4_lut (.I0(n4551[247]), .I1(n1186), .I2(n22943), 
            .I3(n9513), .O(n12185));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8075_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8074_3_lut_4_lut (.I0(n4551[246]), .I1(n1187), .I2(n22943), 
            .I3(n9513), .O(n12184));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8074_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_553_i8_3_lut (.I0(n4551[135]), .I1(n4551[151]), .I2(address_c_0), 
            .I3(GND_net), .O(n4098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_553_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8073_3_lut_4_lut (.I0(n4551[245]), .I1(n1188), .I2(n22943), 
            .I3(n9513), .O(n12183));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8073_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8072_3_lut_4_lut (.I0(n4551[244]), .I1(n1189), .I2(n22943), 
            .I3(n9513), .O(n12182));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8072_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8071_3_lut_4_lut (.I0(n4551[243]), .I1(n1190), .I2(n22943), 
            .I3(n9513), .O(n12181));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8071_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8070_3_lut_4_lut (.I0(n4551[242]), .I1(n1191), .I2(n22943), 
            .I3(n9513), .O(n12180));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8070_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8069_3_lut_4_lut (.I0(n4551[241]), .I1(n1192), .I2(n22943), 
            .I3(n9513), .O(n12179));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8069_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8068_3_lut_4_lut (.I0(n4551[240]), .I1(n1193), .I2(n22943), 
            .I3(n9513), .O(n12178));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8068_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8067_3_lut_4_lut (.I0(n4551[239]), .I1(n1194), .I2(n22943), 
            .I3(n9513), .O(n12177));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8067_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8066_3_lut_4_lut (.I0(n4551[238]), .I1(n1195), .I2(n22943), 
            .I3(n9513), .O(n12176));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8066_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8065_3_lut_4_lut (.I0(n4551[237]), .I1(n1196), .I2(n22943), 
            .I3(n9513), .O(n12175));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8065_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8064_3_lut_4_lut (.I0(n4551[236]), .I1(n1197), .I2(n22943), 
            .I3(n9513), .O(n12174));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8064_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8063_3_lut_4_lut (.I0(n4551[235]), .I1(n1198), .I2(n22943), 
            .I3(n9513), .O(n12173));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8063_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8062_3_lut_4_lut (.I0(n4551[234]), .I1(n1199), .I2(n22943), 
            .I3(n9513), .O(n12172));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8062_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8061_3_lut_4_lut (.I0(n4551[233]), .I1(n1200), .I2(n22943), 
            .I3(n9513), .O(n12171));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8061_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8060_3_lut_4_lut (.I0(n4551[232]), .I1(n1201), .I2(n22943), 
            .I3(n9513), .O(n12170));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8060_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20298_2_lut (.I0(\ootx_crc32_o[0] [15]), .I1(address_c_0), 
            .I2(GND_net), .I3(GND_net), .O(n24666));
    defparam i20298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8059_3_lut_4_lut (.I0(n4551[231]), .I1(n1202), .I2(n22943), 
            .I3(n9513), .O(n12169));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8059_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8058_3_lut_4_lut (.I0(n4551[230]), .I1(n1203), .I2(n22943), 
            .I3(n9513), .O(n12168));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8058_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 n25201_bdd_4_lut (.I0(n25201), .I1(n24233), .I2(n3729), .I3(address_c_4), 
            .O(n25204));
    defparam n25201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8057_3_lut_4_lut (.I0(n4551[229]), .I1(n1204), .I2(n22943), 
            .I3(n9513), .O(n12167));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8057_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8056_3_lut_4_lut (.I0(n4551[228]), .I1(n1205), .I2(n22943), 
            .I3(n9513), .O(n12166));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8056_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_475_i16_3_lut (.I0(n4568[15]), .I1(n4568[31]), .I2(address_c_0), 
            .I3(GND_net), .O(n3093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_561_i16_3_lut (.I0(n4568[95]), .I1(n4568[111]), .I2(address_c_0), 
            .I3(GND_net), .O(n4218));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8055_3_lut_4_lut (.I0(n4551[227]), .I1(n1206), .I2(n22943), 
            .I3(n9513), .O(n12165));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8055_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8054_3_lut_4_lut (.I0(n4551[226]), .I1(n1207), .I2(n22943), 
            .I3(n9513), .O(n12164));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8054_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8053_3_lut_4_lut (.I0(n4551[225]), .I1(n1208), .I2(n22943), 
            .I3(n9513), .O(n12163));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8053_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8052_3_lut_4_lut (.I0(n4551[224]), .I1(n1209), .I2(n22943), 
            .I3(n9513), .O(n12162));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8052_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_563_i16_3_lut (.I0(n4568[63]), .I1(n4568[79]), .I2(address_c_0), 
            .I3(GND_net), .O(n4237));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8051_3_lut_4_lut (.I0(n4551[223]), .I1(n1210), .I2(n22943), 
            .I3(n9513), .O(n12161));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8051_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8050_3_lut_4_lut (.I0(n4551[222]), .I1(n1211), .I2(n22943), 
            .I3(n9513), .O(n12160));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8050_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8049_3_lut_4_lut (.I0(n4551[221]), .I1(n1212), .I2(n22943), 
            .I3(n9513), .O(n12159));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8049_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20297_2_lut (.I0(\ootx_crc32_o[0] [14]), .I1(address_c_0), 
            .I2(GND_net), .I3(GND_net), .O(n24665));
    defparam i20297_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8048_3_lut_4_lut (.I0(n4551[220]), .I1(n1213), .I2(n22943), 
            .I3(n9513), .O(n12158));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8048_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8047_3_lut_4_lut (.I0(n4551[219]), .I1(n1214), .I2(n22943), 
            .I3(n9513), .O(n12157));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8047_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8046_3_lut_4_lut (.I0(n4551[218]), .I1(n1215), .I2(n22943), 
            .I3(n9513), .O(n12156));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8046_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8045_3_lut_4_lut (.I0(n4551[217]), .I1(n1216), .I2(n22943), 
            .I3(n9513), .O(n12155));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8045_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8044_3_lut_4_lut (.I0(n4551[216]), .I1(n1217), .I2(n22943), 
            .I3(n9513), .O(n12154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8044_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8043_3_lut_4_lut (.I0(n4551[215]), .I1(n1218), .I2(n22943), 
            .I3(n9513), .O(n12153));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8043_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8042_3_lut_4_lut (.I0(n4551[214]), .I1(n1219), .I2(n22943), 
            .I3(n9513), .O(n12152));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8042_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8041_3_lut_4_lut (.I0(n4551[213]), .I1(n1220), .I2(n22943), 
            .I3(n9513), .O(n12151));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8041_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8040_3_lut_4_lut (.I0(n4551[212]), .I1(n1221), .I2(n22943), 
            .I3(n9513), .O(n12150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8040_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8039_3_lut_4_lut (.I0(n4551[211]), .I1(n1222), .I2(n22943), 
            .I3(n9513), .O(n12149));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8039_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8038_3_lut_4_lut (.I0(n4551[210]), .I1(n1223), .I2(n22943), 
            .I3(n9513), .O(n12148));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8038_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8037_3_lut_4_lut (.I0(n4551[209]), .I1(n1224), .I2(n22943), 
            .I3(n9513), .O(n12147));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8037_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8036_3_lut_4_lut (.I0(n4551[208]), .I1(n1225), .I2(n22943), 
            .I3(n9513), .O(n12146));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8036_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_475_i15_3_lut (.I0(n4568[14]), .I1(n4568[30]), .I2(address_c_0), 
            .I3(GND_net), .O(n3094));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8035_3_lut_4_lut (.I0(n4551[207]), .I1(n1226), .I2(n22943), 
            .I3(n9513), .O(n12145));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8035_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8034_3_lut_4_lut (.I0(n4551[206]), .I1(n1227), .I2(n22943), 
            .I3(n9513), .O(n12144));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8034_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8033_3_lut_4_lut (.I0(n4551[205]), .I1(n1228), .I2(n22943), 
            .I3(n9513), .O(n12143));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8033_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_561_i15_3_lut (.I0(n4568[94]), .I1(n4568[110]), .I2(address_c_0), 
            .I3(GND_net), .O(n4219));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8032_3_lut_4_lut (.I0(n4551[204]), .I1(n1229), .I2(n22943), 
            .I3(n9513), .O(n12142));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8032_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8031_3_lut_4_lut (.I0(n4551[203]), .I1(n1230), .I2(n22943), 
            .I3(n9513), .O(n12141));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8031_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8030_3_lut_4_lut (.I0(n4551[202]), .I1(n1231), .I2(n22943), 
            .I3(n9513), .O(n12140));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8030_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8029_3_lut_4_lut (.I0(n4551[201]), .I1(n1232), .I2(n22943), 
            .I3(n9513), .O(n12139));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8029_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8028_3_lut_4_lut (.I0(n4551[200]), .I1(n1233), .I2(n22943), 
            .I3(n9513), .O(n12138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8028_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8027_3_lut_4_lut (.I0(n4551[199]), .I1(n1234), .I2(n22943), 
            .I3(n9513), .O(n12137));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8027_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_563_i15_3_lut (.I0(n4568[62]), .I1(n4568[78]), .I2(address_c_0), 
            .I3(GND_net), .O(n4238));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20296_2_lut (.I0(\ootx_crc32_o[0] [13]), .I1(address_c_0), 
            .I2(GND_net), .I3(GND_net), .O(n24664));
    defparam i20296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8026_3_lut_4_lut (.I0(n4551[198]), .I1(n1235), .I2(n22943), 
            .I3(n9513), .O(n12136));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8026_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8025_3_lut_4_lut (.I0(n4551[197]), .I1(n1236), .I2(n22943), 
            .I3(n9513), .O(n12135));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8025_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8024_3_lut_4_lut (.I0(n4551[196]), .I1(n1237), .I2(n22943), 
            .I3(n9513), .O(n12134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8024_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8023_3_lut_4_lut (.I0(n4551[195]), .I1(n1238), .I2(n22943), 
            .I3(n9513), .O(n12133));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8023_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8022_3_lut_4_lut (.I0(n4551[194]), .I1(n1239), .I2(n22943), 
            .I3(n9513), .O(n12132));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8022_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8021_3_lut_4_lut (.I0(n4551[193]), .I1(n1240), .I2(n22943), 
            .I3(n9513), .O(n12131));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8021_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8020_3_lut_4_lut (.I0(n4551[192]), .I1(n1241), .I2(n22943), 
            .I3(n9513), .O(n12130));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8020_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8019_3_lut_4_lut (.I0(n4551[191]), .I1(n1242), .I2(n22943), 
            .I3(n9513), .O(n12129));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8019_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_475_i14_3_lut (.I0(n4568[13]), .I1(n4568[29]), .I2(address_c_0), 
            .I3(GND_net), .O(n3095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8018_3_lut_4_lut (.I0(n4551[190]), .I1(n1243), .I2(n22943), 
            .I3(n9513), .O(n12128));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8018_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8017_3_lut_4_lut (.I0(n4551[189]), .I1(n1244), .I2(n22943), 
            .I3(n9513), .O(n12127));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8017_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8016_3_lut_4_lut (.I0(n4551[188]), .I1(n1245), .I2(n22943), 
            .I3(n9513), .O(n12126));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8016_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8015_3_lut_4_lut (.I0(n4551[187]), .I1(n1246), .I2(n22943), 
            .I3(n9513), .O(n12125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8015_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8014_3_lut_4_lut (.I0(n4551[186]), .I1(n1247), .I2(n22943), 
            .I3(n9513), .O(n12124));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8014_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8013_3_lut_4_lut (.I0(n4551[185]), .I1(n1248), .I2(n22943), 
            .I3(n9513), .O(n12123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8013_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8012_3_lut_4_lut (.I0(n4551[184]), .I1(n1249), .I2(n22943), 
            .I3(n9513), .O(n12122));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8012_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8011_3_lut_4_lut (.I0(n4551[183]), .I1(n1250), .I2(n22943), 
            .I3(n9513), .O(n12121));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8011_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8010_3_lut_4_lut (.I0(n4551[182]), .I1(n1251), .I2(n22943), 
            .I3(n9513), .O(n12120));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8010_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8009_3_lut_4_lut (.I0(n4551[181]), .I1(n1252), .I2(n22943), 
            .I3(n9513), .O(n12119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8009_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_561_i14_3_lut (.I0(n4568[93]), .I1(n4568[109]), .I2(address_c_0), 
            .I3(GND_net), .O(n4220));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_561_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8008_3_lut_4_lut (.I0(n4551[180]), .I1(n1253), .I2(n22943), 
            .I3(n9513), .O(n12118));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8008_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8007_3_lut_4_lut (.I0(n4551[179]), .I1(n1254), .I2(n22943), 
            .I3(n9513), .O(n12117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8007_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8006_3_lut_4_lut (.I0(n4551[178]), .I1(n1255), .I2(n22943), 
            .I3(n9513), .O(n12116));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8006_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_563_i14_3_lut (.I0(n4568[61]), .I1(n4568[77]), .I2(address_c_0), 
            .I3(GND_net), .O(n4239));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_563_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14599_3_lut_4_lut (.I0(n4551[177]), .I1(n1256), .I2(n22943), 
            .I3(n9513), .O(n12115));
    defparam i14599_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i20295_2_lut (.I0(\ootx_crc32_o[0] [12]), .I1(address_c_0), 
            .I2(GND_net), .I3(GND_net), .O(n24663));
    defparam i20295_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8004_3_lut_4_lut (.I0(n4551[176]), .I1(n1257), .I2(n22943), 
            .I3(n9513), .O(n12114));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8004_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i8003_3_lut_4_lut (.I0(n4551[175]), .I1(n1258), .I2(n22943), 
            .I3(n9513), .O(n12113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8003_3_lut_4_lut.LUT_INIT = 16'hacaa;
    GND i1 (.Y(GND_net));
    SB_LUT4 i8002_3_lut_4_lut (.I0(n4551[174]), .I1(n1259), .I2(n22943), 
            .I3(n9513), .O(n12112));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8002_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_475_i13_3_lut (.I0(n4568[12]), .I1(n4568[28]), .I2(address_c_0), 
            .I3(GND_net), .O(n3096));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(59[2] 95[15])
    defparam mux_475_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8001_3_lut_4_lut (.I0(n4551[173]), .I1(n1260), .I2(n22943), 
            .I3(n9513), .O(n12111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    defparam i8001_3_lut_4_lut.LUT_INIT = 16'hacaa;
    
endmodule
//
// Verilog Description of module lighthouse_ootx_decoder_default
//

module lighthouse_ootx_decoder_default (\lighthouse[0] , n6333, counter_from_last_rise, 
            GND_net, \ootx_payload_o[1][0] , clock_c, n1, n1_adj_1, 
            n1000, data, n1194, \ootx_payloads_N_1730[1] , n2851, 
            bit_counters_0_7, bit_counters_1_7, bit_counters_0_8, bit_counters_1_8, 
            bit_counters_0_9, bit_counters_1_9, \ootx_payloads_N_1730[2] , 
            n24018, \ootx_payloads_N_1699[4] , n13221, reset_c, new_data, 
            ootx_payloads_N_1744, bit_counters_0_10, bit_counters_1_10, 
            \ootx_payloads_N_1730[3] , n337, n998, n1195, n996, n1196, 
            n994, n1197, VCC_net, n992, n1198, n766, n1311, n13, 
            n990, n1199, n988, n1200, n1_adj_2, n9797, n23974, 
            n8, bit_counters_0_19, bit_counters_1_19, n23003, data_counters_0_0, 
            n23005, data_counters_0_1, n23007, data_counters_0_2, n23009, 
            data_counters_0_3, n23011, data_counters_0_4, n23013, data_counters_0_5, 
            n23015, data_counters_0_6, n23017, data_counters_0_7, n23019, 
            data_counters_0_8, n23021, data_counters_0_9, n23023, data_counters_0_10, 
            n1_adj_3, n23025, data_counters_0_11, n23027, data_counters_0_12, 
            n23029, data_counters_0_13, n23031, data_counters_0_14, 
            n23033, data_counters_0_15, n23035, data_counters_0_16, 
            n23037, data_counters_0_17, n23039, data_counters_0_18, 
            n23041, data_counters_0_19, n23043, data_counters_0_20, 
            n23045, data_counters_0_21, n23047, data_counters_0_22, 
            n23049, data_counters_0_23, n23051, data_counters_0_24, 
            n23053, data_counters_0_25, n23055, data_counters_0_26, 
            n23057, data_counters_0_27, n23059, data_counters_0_28, 
            n23061, data_counters_0_29, n23063, data_counters_0_30, 
            n23065, data_counters_1_0, n23067, data_counters_1_1, n23069, 
            data_counters_1_2, n23071, data_counters_1_3, n23073, data_counters_1_4, 
            n23075, data_counters_1_5, n23077, data_counters_1_6, n23079, 
            data_counters_1_7, n23081, data_counters_1_8, n23083, data_counters_1_9, 
            n23085, data_counters_1_10, n23087, data_counters_1_11, 
            n23089, data_counters_1_12, n23091, data_counters_1_13, 
            n23093, data_counters_1_14, n23095, data_counters_1_15, 
            n23097, data_counters_1_16, n23099, data_counters_1_17, 
            n23101, data_counters_1_18, n23103, data_counters_1_19, 
            n23105, data_counters_1_20, n23107, data_counters_1_21, 
            n23109, data_counters_1_22, n23111, data_counters_1_23, 
            n23113, data_counters_1_24, n23115, data_counters_1_25, 
            n23117, data_counters_1_26, n23119, data_counters_1_27, 
            n23121, data_counters_1_28, n23123, data_counters_1_29, 
            n23125, data_counters_1_30, n23475, bit_counters_0_0, n23477, 
            bit_counters_0_1, n23479, bit_counters_0_2, n23481, bit_counters_0_3, 
            n23483, bit_counters_0_4, n23485, bit_counters_0_5, n23487, 
            bit_counters_0_6, n23489, n23491, n23493, n23495, n23497, 
            bit_counters_0_11, n23499, bit_counters_0_12, n23501, bit_counters_0_13, 
            n23503, bit_counters_0_14, n23505, bit_counters_0_15, n23507, 
            bit_counters_0_16, n23509, bit_counters_0_17, n23469, bit_counters_0_18, 
            n23463, n23457, bit_counters_0_20, n23451, bit_counters_0_21, 
            n23445, bit_counters_0_22, n23439, bit_counters_0_23, n23433, 
            bit_counters_0_24, n23427, bit_counters_0_25, n23421, bit_counters_0_26, 
            n23415, bit_counters_0_27, n23409, bit_counters_0_28, n23399, 
            bit_counters_0_29, n23389, bit_counters_0_30, n23511, bit_counters_1_0, 
            n23513, bit_counters_1_1, n23515, bit_counters_1_2, n23517, 
            bit_counters_1_3, n23519, bit_counters_1_4, n23521, bit_counters_1_5, 
            n23523, bit_counters_1_6, n23525, n23527, n23529, n23531, 
            n23533, bit_counters_1_11, n23535, bit_counters_1_12, n23537, 
            bit_counters_1_13, n23539, bit_counters_1_14, n23541, bit_counters_1_15, 
            n23543, bit_counters_1_16, n23545, bit_counters_1_17, n23471, 
            bit_counters_1_18, n23465, n23459, bit_counters_1_20, n23453, 
            bit_counters_1_21, n23447, bit_counters_1_22, n23441, bit_counters_1_23, 
            n23435, bit_counters_1_24, n23429, bit_counters_1_25, n23423, 
            bit_counters_1_26, n23417, bit_counters_1_27, n986, n1201, 
            n35, n23411, bit_counters_1_28, n23401, bit_counters_1_29, 
            n23391, bit_counters_1_30, n23697, n23639, payload_lengths_0_0, 
            n23641, payload_lengths_1_0, n8_adj_4, n8_adj_5, n8_adj_6, 
            n2282, n8_adj_7, n984, n1202, n8_adj_8, \counter_from_last_rise[6] , 
            n8_adj_9, \counter_from_last_rise[7] , n8_adj_10, \counter_from_last_rise[8] , 
            n8_adj_11, \counter_from_last_rise[9] , n8_adj_12, \counter_from_last_rise[10] , 
            n8_adj_13, \counter_from_last_rise[11] , n8_adj_14, \counter_from_last_rise[12] , 
            n8_adj_15, n8_adj_16, n8_adj_17, n8_adj_18, n8_adj_19, 
            n8_adj_20, n8_adj_21, \counter_from_last_rise[19] , n8_adj_22, 
            \counter_from_last_rise[20] , n8_adj_23, \counter_from_last_rise[21] , 
            n8_adj_24, \counter_from_last_rise[22] , n8_adj_25, \counter_from_last_rise[23] , 
            n8_adj_26, \counter_from_last_rise[24] , n8_adj_27, \counter_from_last_rise[25] , 
            n8_adj_28, \counter_from_last_rise[26] , n8_adj_29, \counter_from_last_rise[27] , 
            n8_adj_30, \counter_from_last_rise[28] , n8_adj_31, \counter_from_last_rise[29] , 
            n23407, \counter_from_last_rise[30] , n23397, \counter_from_last_rise[31] , 
            n12201, \ootx_payload_o[0][263] , n12200, \ootx_payload_o[0][262] , 
            n12199, \ootx_payload_o[0][261] , n12198, \ootx_payload_o[0][260] , 
            n12197, \ootx_payload_o[0][259] , n12196, \ootx_payload_o[0][258] , 
            n12195, \ootx_payload_o[0][257] , n12194, \ootx_payload_o[0][256] , 
            n12193, \ootx_payload_o[0][255] , n12192, \ootx_payload_o[0][254] , 
            n12191, \ootx_payload_o[0][253] , n12190, \ootx_payload_o[0][252] , 
            n12189, \ootx_payload_o[0][251] , n12188, \ootx_payload_o[0][250] , 
            n12187, \ootx_payload_o[0][249] , n12186, \ootx_payload_o[0][248] , 
            n12185, \ootx_payload_o[0][247] , n12184, \ootx_payload_o[0][246] , 
            n12183, \ootx_payload_o[0][245] , n12182, \ootx_payload_o[0][244] , 
            n12181, \ootx_payload_o[0][243] , n12180, \ootx_payload_o[0][242] , 
            n12179, \ootx_payload_o[0][241] , n12178, \ootx_payload_o[0][240] , 
            n12177, \ootx_payload_o[0][239] , n12176, \ootx_payload_o[0][238] , 
            n12175, \ootx_payload_o[0][237] , n12174, \ootx_payload_o[0][236] , 
            n12173, \ootx_payload_o[0][235] , n12172, \ootx_payload_o[0][234] , 
            n12171, \ootx_payload_o[0][233] , n12170, \ootx_payload_o[0][232] , 
            n12169, \ootx_payload_o[0][231] , n12168, \ootx_payload_o[0][230] , 
            n12167, \ootx_payload_o[0][229] , n12166, \ootx_payload_o[0][228] , 
            n12165, \ootx_payload_o[0][227] , n12164, \ootx_payload_o[0][226] , 
            n12163, \ootx_payload_o[0][225] , n12162, \ootx_payload_o[0][224] , 
            n12161, \ootx_payload_o[0][223] , n12160, \ootx_payload_o[0][222] , 
            n12159, \ootx_payload_o[0][221] , n12158, \ootx_payload_o[0][220] , 
            n12157, \ootx_payload_o[0][219] , n12156, \ootx_payload_o[0][218] , 
            n12155, \ootx_payload_o[0][217] , n12154, \ootx_payload_o[0][216] , 
            n12153, \ootx_payload_o[0][215] , n12152, \ootx_payload_o[0][214] , 
            n12151, \ootx_payload_o[0][213] , n12150, \ootx_payload_o[0][212] , 
            n12149, \ootx_payload_o[0][211] , n12148, \ootx_payload_o[0][210] , 
            n12147, \ootx_payload_o[0][209] , n12146, \ootx_payload_o[0][208] , 
            n12145, \ootx_payload_o[0][207] , n12144, \ootx_payload_o[0][206] , 
            n12143, \ootx_payload_o[0][205] , n12142, \ootx_payload_o[0][204] , 
            n12141, \ootx_payload_o[0][203] , n12140, \ootx_payload_o[0][202] , 
            n12139, \ootx_payload_o[0][201] , n12138, \ootx_payload_o[0][200] , 
            n12137, \ootx_payload_o[0][199] , n12136, \ootx_payload_o[0][198] , 
            n12135, \ootx_payload_o[0][197] , n12134, \ootx_payload_o[0][196] , 
            n12133, \ootx_payload_o[0][195] , n12132, \ootx_payload_o[0][194] , 
            n12131, \ootx_payload_o[0][193] , n12130, \ootx_payload_o[0][192] , 
            n12129, \ootx_payload_o[0][191] , n12128, \ootx_payload_o[0][190] , 
            n12127, \ootx_payload_o[0][189] , n12126, \ootx_payload_o[0][188] , 
            n12125, \ootx_payload_o[0][187] , n12124, \ootx_payload_o[0][186] , 
            n12123, \ootx_payload_o[0][185] , n12122, \ootx_payload_o[0][184] , 
            n12121, \ootx_payload_o[0][183] , n12120, \ootx_payload_o[0][182] , 
            n12119, \ootx_payload_o[0][181] , n12118, \ootx_payload_o[0][180] , 
            n12117, \ootx_payload_o[0][179] , n12116, \ootx_payload_o[0][178] , 
            n12115, \ootx_payload_o[0][177] , n12114, \ootx_payload_o[0][176] , 
            n12113, \ootx_payload_o[0][175] , n12112, \ootx_payload_o[0][174] , 
            n12111, \ootx_payload_o[0][173] , n12110, \ootx_payload_o[0][172] , 
            n12109, \ootx_payload_o[0][171] , n12108, \ootx_payload_o[0][170] , 
            n12107, \ootx_payload_o[0][169] , n12106, \ootx_payload_o[0][168] , 
            n12105, \ootx_payload_o[0][167] , n12104, \ootx_payload_o[0][166] , 
            n12103, \ootx_payload_o[0][165] , n12102, \ootx_payload_o[0][164] , 
            n12101, \ootx_payload_o[0][163] , n12100, \ootx_payload_o[0][162] , 
            n12099, \ootx_payload_o[0][161] , n12098, \ootx_payload_o[0][160] , 
            n12097, \ootx_payload_o[0][159] , n12096, \ootx_payload_o[0][158] , 
            n12095, \ootx_payload_o[0][157] , n12094, \ootx_payload_o[0][156] , 
            n12093, \ootx_payload_o[0][155] , n12092, \ootx_payload_o[0][154] , 
            n12091, \ootx_payload_o[0][153] , n12090, \ootx_payload_o[0][152] , 
            n12089, \ootx_payload_o[0][151] , n12088, \ootx_payload_o[0][150] , 
            n12087, \ootx_payload_o[0][149] , n12086, \ootx_payload_o[0][148] , 
            n12085, \ootx_payload_o[0][147] , n12084, \ootx_payload_o[0][146] , 
            n12083, \ootx_payload_o[0][145] , n12082, \ootx_payload_o[0][144] , 
            n12081, \ootx_payload_o[0][143] , n12080, \ootx_payload_o[0][142] , 
            n12079, \ootx_payload_o[0][141] , n12078, \ootx_payload_o[0][140] , 
            n12077, \ootx_payload_o[0][139] , n12076, \ootx_payload_o[0][138] , 
            n12075, \ootx_payload_o[0][137] , n12074, \ootx_payload_o[0][136] , 
            n12073, \ootx_payload_o[0][135] , n12072, \ootx_payload_o[0][134] , 
            n12071, \ootx_payload_o[0][133] , n12070, \ootx_payload_o[0][132] , 
            n12069, \ootx_payload_o[0][131] , n12068, \ootx_payload_o[0][130] , 
            n12067, \ootx_payload_o[0][129] , n12066, \ootx_payload_o[0][128] , 
            n12065, \ootx_payload_o[0][127] , n12064, \ootx_payload_o[0][126] , 
            n12063, \ootx_payload_o[0][125] , n12062, \ootx_payload_o[0][124] , 
            n12061, \ootx_payload_o[0][123] , n12060, \ootx_payload_o[0][122] , 
            n12059, \ootx_payload_o[0][121] , n12058, \ootx_payload_o[0][120] , 
            n12057, \ootx_payload_o[0][119] , n12056, \ootx_payload_o[0][118] , 
            n12055, \ootx_payload_o[0][117] , n12054, \ootx_payload_o[0][116] , 
            n12053, \ootx_payload_o[0][115] , n12052, \ootx_payload_o[0][114] , 
            n12051, \ootx_payload_o[0][113] , n12050, \ootx_payload_o[0][112] , 
            n12049, \ootx_payload_o[0][111] , n12048, \ootx_payload_o[0][110] , 
            n12047, \ootx_payload_o[0][109] , n12046, \ootx_payload_o[0][108] , 
            n12045, \ootx_payload_o[0][107] , n12044, \ootx_payload_o[0][106] , 
            n12043, \ootx_payload_o[0][105] , n12042, \ootx_payload_o[0][104] , 
            n12041, \ootx_payload_o[0][103] , n12040, \ootx_payload_o[0][102] , 
            n12039, \ootx_payload_o[0][101] , n12038, \ootx_payload_o[0][100] , 
            n12037, \ootx_payload_o[0][99] , n12036, \ootx_payload_o[0][98] , 
            n12035, \ootx_payload_o[0][97] , n12034, \ootx_payload_o[0][96] , 
            n12033, \ootx_payload_o[0][95] , n12032, \ootx_payload_o[0][94] , 
            n12031, \ootx_payload_o[0][93] , n12030, \ootx_payload_o[0][92] , 
            n12029, \ootx_payload_o[0][91] , n12028, \ootx_payload_o[0][90] , 
            n12027, \ootx_payload_o[0][89] , n12026, \ootx_payload_o[0][88] , 
            n12025, \ootx_payload_o[0][87] , n12024, \ootx_payload_o[0][86] , 
            n12023, \ootx_payload_o[0][85] , n12022, \ootx_payload_o[0][84] , 
            n12021, \ootx_payload_o[0][83] , n12020, \ootx_payload_o[0][82] , 
            n12019, \ootx_payload_o[0][81] , n12018, \ootx_payload_o[0][80] , 
            n12017, \ootx_payload_o[0][79] , n12016, \ootx_payload_o[0][78] , 
            n12015, \ootx_payload_o[0][77] , n12014, \ootx_payload_o[0][76] , 
            n12013, \ootx_payload_o[0][75] , n12012, \ootx_payload_o[0][74] , 
            n12011, \ootx_payload_o[0][73] , n12010, \ootx_payload_o[0][72] , 
            n12009, \ootx_payload_o[0][71] , n12008, \ootx_payload_o[0][70] , 
            n12007, \ootx_payload_o[0][69] , n12006, \ootx_payload_o[0][68] , 
            n12005, \ootx_payload_o[0][67] , n12004, \ootx_payload_o[0][66] , 
            n12003, \ootx_payload_o[0][65] , n12002, \ootx_payload_o[0][64] , 
            n12001, \ootx_payload_o[0][63] , n12000, \ootx_payload_o[0][62] , 
            n11999, \ootx_payload_o[0][61] , n11998, \ootx_payload_o[0][60] , 
            n11997, \ootx_payload_o[0][59] , n11996, \ootx_payload_o[0][58] , 
            n11995, \ootx_payload_o[0][57] , n11994, \ootx_payload_o[0][56] , 
            n11993, \ootx_payload_o[0][55] , n11992, \ootx_payload_o[0][54] , 
            n11991, \ootx_payload_o[0][53] , n11990, \ootx_payload_o[0][52] , 
            n938, n1225, n11989, \ootx_payload_o[0][51] , n11988, 
            \ootx_payload_o[0][50] , n11987, \ootx_payload_o[0][49] , 
            n11986, \ootx_payload_o[0][48] , n11985, \ootx_payload_o[0][47] , 
            n11984, \ootx_payload_o[0][46] , n11983, \ootx_payload_o[0][45] , 
            n958, n1215, n11982, \ootx_payload_o[0][44] , n30, n11981, 
            \ootx_payload_o[0][43] , n11980, \ootx_payload_o[0][42] , 
            n11979, \ootx_payload_o[0][41] , n11978, \ootx_payload_o[0][40] , 
            n11977, \ootx_payload_o[0][39] , n982, n1203, n11976, 
            \ootx_payload_o[0][38] , n11975, \ootx_payload_o[0][37] , 
            n11974, \ootx_payload_o[0][36] , n11973, \ootx_payload_o[0][35] , 
            sensor_state, n11972, \ootx_payload_o[0][34] , n11971, \ootx_payload_o[0][33] , 
            n11970, \ootx_payload_o[0][32] , n11969, \ootx_payload_o[0][31] , 
            n11968, \ootx_payload_o[0][30] , n11967, \ootx_payload_o[0][29] , 
            n11966, \ootx_payload_o[0][28] , n11965, \ootx_payload_o[0][27] , 
            n11964, \ootx_payload_o[0][26] , n11963, \ootx_payload_o[0][25] , 
            n11962, \ootx_payload_o[0][24] , n11961, \ootx_payload_o[0][23] , 
            n11960, \ootx_payload_o[0][22] , n11959, \ootx_payload_o[0][21] , 
            n680, n1354, n712, n1338, \ootx_payloads_N_1699[5] , \ootx_payloads_N_1699[3] , 
            \ootx_payloads_N_1699[15] , n34, n11958, \ootx_payload_o[0][20] , 
            n11957, \ootx_payload_o[0][19] , n11956, \ootx_payload_o[0][18] , 
            n11955, \ootx_payload_o[0][17] , n11954, \ootx_payload_o[0][16] , 
            n11953, \ootx_payload_o[0][15] , n11952, \ootx_payload_o[0][14] , 
            n11951, \ootx_payload_o[0][13] , n11950, \ootx_payload_o[0][12] , 
            n11949, \ootx_payload_o[0][11] , n11948, \ootx_payload_o[0][10] , 
            n11947, \ootx_payload_o[0][9] , n11946, \ootx_payload_o[0][8] , 
            n11945, \ootx_payload_o[0][7] , n11944, \ootx_payload_o[0][6] , 
            n11943, \ootx_payload_o[0][5] , n11942, \ootx_payload_o[0][4] , 
            n11941, \ootx_payload_o[0][3] , n11940, \ootx_payload_o[0][2] , 
            n11939, \ootx_payload_o[0][1] , \ootx_crc32_o[1] , \ootx_crc32_o[0] , 
            n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
            n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
            n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
            n640, n1374, n724, n928, n1230, n1204, n1205, n1206, 
            n1207, n1208, n1209, n1210, n1332, n1211, n1212, n1213, 
            \ootx_payloads_N_1699[6] , \ootx_payloads_N_1699[7] , \ootx_payloads_N_1699[8] , 
            n1010, n1214, n754, n764, n672, \ootx_states[0] , n638, 
            n1375, ootx_payloads_1_263, n926, n1231, n670, n1312, 
            n20, ootx_payloads_1_262, n924, n1232, n636, n1376, 
            n668, n922, n1233, n634, n1377, n666, n920, n1234, 
            n632, n1378, n664, n918, n1235, n662, n916, n1236, 
            n752, n1318, n660, n914, n1237, n658, n678, n1355, 
            n912, n1238, n630, n1379, ootx_payloads_1_261, ootx_payloads_1_260, 
            n656, ootx_payloads_1_259, n910, n1239, n654, n1008, 
            n676, n1356, n908, n1240, ootx_payloads_1_258, ootx_payloads_1_257, 
            ootx_payloads_1_256, n628, n1380, ootx_payloads_1_255, \ootx_payloads_N_1699[30] , 
            n9200, \ootx_payloads_N_1699[9] , \ootx_payloads_N_1699[13] , 
            \ootx_payloads_N_1699[12] , \ootx_payloads_N_1699[11] , ootx_payloads_1_254, 
            ootx_payloads_1_253, ootx_payloads_1_252, ootx_payloads_1_251, 
            n652, n906, n1241, ootx_payloads_1_250, ootx_payloads_1_249, 
            \ootx_payloads_N_1699[10] , \ootx_payloads_N_1699[14] , n650, 
            n626, n1381, n904, n1242, n648, n980, n624, n1382, 
            ootx_payloads_1_248, ootx_payloads_1_247, n902, n1243, n900, 
            n1244, n978, n674, n1357, n19, n622, n1383, ootx_payloads_1_246, 
            ootx_payloads_1_245, n898, n1245, ootx_payloads_1_244, n896, 
            n1246, n620, n1384, n6355, n894, n1247, n6356, n6357, 
            \ootx_payloads_N_1730[4] , n6358, n750, n1319, n618, n1385, 
            n892, n1248, n6359, ootx_payloads_1_243, n6361, n890, 
            n1249, ootx_payloads_1_242, n6362, n616, n1386, ootx_payloads_1_241, 
            ootx_payloads_1_240, ootx_payloads_1_239, n1006, n888, n1250, 
            ootx_payloads_1_238, ootx_payloads_1_237, n886, n1251, n614, 
            n1387, n22943, n976, ootx_payloads_1_236, n884, n1252, 
            ootx_payloads_1_235, n882, n1253, ootx_payloads_1_234, n1358, 
            n612, n1388, n880, n1254, n748, n1320, n974, n878, 
            n1255, n1004, n13329, data_N_1808, n6363, n6364, n6365, 
            ootx_payloads_1_233, sensor_N_132, n876, n1256, ootx_payloads_1_232, 
            n610, n1389, ootx_payloads_1_231, n874, n1257, n872, 
            n1258, n608, n1390, n870, n1259, n746, n1321, n606, 
            n1391, n604, n1392, n710, n1339, n966, n868, n1260, 
            n602, n1393, n744, n1322, n866, n1261, n600, n1394, 
            n864, n1262, n598, n1395, ootx_payloads_1_230, ootx_payloads_1_229, 
            ootx_payloads_1_228, ootx_payloads_1_227, n596, n1396, n594, 
            n1397, ootx_payloads_1_226, ootx_payloads_1_225, ootx_payloads_1_224, 
            n592, n1398, ootx_payloads_1_223, n742, n1323, n862, 
            n1263, n590, n1399, ootx_payloads_1_222, ootx_payloads_1_221, 
            \ootx_payload_o[1][1] , ootx_payloads_1_220, ootx_payloads_1_219, 
            ootx_payloads_1_218, n588, n1400, ootx_payloads_1_217, ootx_payloads_1_216, 
            \ootx_payload_o[1][2] , \ootx_payload_o[1][3] , \ootx_payload_o[1][4] , 
            \ootx_payload_o[1][5] , \ootx_payload_o[1][6] , \ootx_payload_o[1][7] , 
            \ootx_payload_o[1][8] , \ootx_payload_o[1][9] , \ootx_payload_o[1][10] , 
            \ootx_payload_o[1][11] , \ootx_payload_o[1][12] , \ootx_payload_o[1][13] , 
            \ootx_payload_o[1][14] , \ootx_payload_o[1][15] , \ootx_payload_o[1][16] , 
            \ootx_payload_o[1][17] , \ootx_payload_o[1][18] , \ootx_payload_o[1][19] , 
            \ootx_payload_o[1][20] , \ootx_payload_o[1][21] , \ootx_payload_o[1][22] , 
            \ootx_payload_o[1][23] , \ootx_payload_o[1][24] , \ootx_payload_o[1][25] , 
            \ootx_payload_o[1][26] , \ootx_payload_o[1][27] , \ootx_payload_o[1][28] , 
            \ootx_payload_o[1][29] , \ootx_payload_o[1][30] , \ootx_payload_o[1][31] , 
            \ootx_payload_o[1][32] , \ootx_payload_o[1][33] , \ootx_payload_o[1][34] , 
            \ootx_payload_o[1][35] , \ootx_payload_o[1][36] , \ootx_payload_o[1][37] , 
            \ootx_payload_o[1][38] , \ootx_payload_o[1][39] , \ootx_payload_o[1][40] , 
            \ootx_payload_o[1][41] , \ootx_payload_o[1][42] , \ootx_payload_o[1][43] , 
            \ootx_payload_o[1][44] , \ootx_payload_o[1][45] , \ootx_payload_o[1][46] , 
            \ootx_payload_o[1][47] , \ootx_payload_o[1][48] , \ootx_payload_o[1][49] , 
            \ootx_payload_o[1][50] , \ootx_payload_o[1][51] , \ootx_payload_o[1][52] , 
            \ootx_payload_o[1][53] , \ootx_payload_o[1][54] , \ootx_payload_o[1][55] , 
            \ootx_payload_o[1][56] , \ootx_payload_o[1][57] , \ootx_payload_o[1][58] , 
            \ootx_payload_o[1][59] , \ootx_payload_o[1][60] , \ootx_payload_o[1][61] , 
            \ootx_payload_o[1][62] , \ootx_payload_o[1][63] , \ootx_payload_o[1][64] , 
            \ootx_payload_o[1][65] , \ootx_payload_o[1][66] , \ootx_payload_o[1][67] , 
            \ootx_payload_o[1][68] , \ootx_payload_o[1][69] , \ootx_payload_o[1][70] , 
            \ootx_payload_o[1][71] , \ootx_payload_o[1][72] , \ootx_payload_o[1][73] , 
            \ootx_payload_o[1][74] , \ootx_payload_o[1][75] , \ootx_payload_o[1][76] , 
            \ootx_payload_o[1][77] , \ootx_payload_o[1][78] , \ootx_payload_o[1][79] , 
            \ootx_payload_o[1][80] , \ootx_payload_o[1][81] , \ootx_payload_o[1][82] , 
            \ootx_payload_o[1][83] , \ootx_payload_o[1][84] , \ootx_payload_o[1][85] , 
            \ootx_payload_o[1][86] , \ootx_payload_o[1][87] , \ootx_payload_o[1][88] , 
            \ootx_payload_o[1][89] , \ootx_payload_o[1][90] , \ootx_payload_o[1][91] , 
            \ootx_payload_o[1][92] , \ootx_payload_o[1][93] , \ootx_payload_o[1][94] , 
            \ootx_payload_o[1][95] , \ootx_payload_o[1][96] , \ootx_payload_o[1][97] , 
            \ootx_payload_o[1][98] , \ootx_payload_o[1][99] , \ootx_payload_o[1][100] , 
            \ootx_payload_o[1][101] , \ootx_payload_o[1][102] , \ootx_payload_o[1][103] , 
            \ootx_payload_o[1][104] , \ootx_payload_o[1][105] , \ootx_payload_o[1][106] , 
            \ootx_payload_o[1][107] , \ootx_payload_o[1][108] , \ootx_payload_o[1][109] , 
            \ootx_payload_o[1][110] , \ootx_payload_o[1][111] , \ootx_payload_o[1][112] , 
            \ootx_payload_o[1][113] , \ootx_payload_o[1][114] , \ootx_payload_o[1][115] , 
            \ootx_payload_o[1][116] , \ootx_payload_o[1][117] , \ootx_payload_o[1][118] , 
            \ootx_payload_o[1][119] , \ootx_payload_o[1][120] , \ootx_payload_o[1][121] , 
            \ootx_payload_o[1][122] , \ootx_payload_o[1][123] , \ootx_payload_o[1][124] , 
            \ootx_payload_o[1][125] , \ootx_payload_o[1][126] , \ootx_payload_o[1][127] , 
            \ootx_payload_o[1][128] , \ootx_payload_o[1][129] , \ootx_payload_o[1][130] , 
            \ootx_payload_o[1][131] , \ootx_payload_o[1][132] , \ootx_payload_o[1][133] , 
            \ootx_payload_o[1][134] , \ootx_payload_o[1][135] , \ootx_payload_o[1][136] , 
            \ootx_payload_o[1][137] , \ootx_payload_o[1][138] , \ootx_payload_o[1][139] , 
            \ootx_payload_o[1][140] , \ootx_payload_o[1][141] , \ootx_payload_o[1][142] , 
            \ootx_payload_o[1][143] , \ootx_payload_o[1][144] , \ootx_payload_o[1][145] , 
            \ootx_payload_o[1][146] , \ootx_payload_o[1][147] , \ootx_payload_o[1][148] , 
            \ootx_payload_o[1][149] , \ootx_payload_o[1][150] , \ootx_payload_o[1][151] , 
            \ootx_payload_o[1][152] , \ootx_payload_o[1][153] , \ootx_payload_o[1][154] , 
            \ootx_payload_o[1][155] , \ootx_payload_o[1][156] , \ootx_payload_o[1][157] , 
            \ootx_payload_o[1][158] , \ootx_payload_o[1][159] , \ootx_payload_o[1][160] , 
            \ootx_payload_o[1][161] , \ootx_payload_o[1][162] , \ootx_payload_o[1][163] , 
            \ootx_payload_o[1][164] , \ootx_payload_o[1][165] , \ootx_payload_o[1][166] , 
            \ootx_payload_o[1][167] , \ootx_payload_o[1][168] , \ootx_payload_o[1][169] , 
            \ootx_payload_o[1][170] , \ootx_payload_o[1][171] , \ootx_payload_o[1][172] , 
            \ootx_payload_o[1][173] , \ootx_payload_o[1][174] , \ootx_payload_o[1][175] , 
            \ootx_payload_o[1][176] , \ootx_payload_o[1][177] , \ootx_payload_o[1][178] , 
            \ootx_payload_o[1][179] , \ootx_payload_o[1][180] , \ootx_payload_o[1][181] , 
            \ootx_payload_o[1][182] , \ootx_payload_o[1][183] , \ootx_payload_o[1][184] , 
            \ootx_payload_o[1][185] , \ootx_payload_o[1][186] , \ootx_payload_o[1][187] , 
            \ootx_payload_o[1][188] , \ootx_payload_o[1][189] , \ootx_payload_o[1][190] , 
            \ootx_payload_o[1][191] , \ootx_payload_o[1][192] , \ootx_payload_o[1][193] , 
            \ootx_payload_o[1][194] , \ootx_payload_o[1][195] , \ootx_payload_o[1][196] , 
            \ootx_payload_o[1][197] , \ootx_payload_o[1][198] , \ootx_payload_o[1][199] , 
            \ootx_payload_o[1][200] , \ootx_payload_o[1][201] , \ootx_payload_o[1][202] , 
            \ootx_payload_o[1][203] , \ootx_payload_o[1][204] , \ootx_payload_o[1][205] , 
            \ootx_payload_o[1][206] , \ootx_payload_o[1][207] , \ootx_payload_o[1][208] , 
            \ootx_payload_o[1][209] , \ootx_payload_o[1][210] , \ootx_payload_o[1][211] , 
            \ootx_payload_o[1][212] , \ootx_payload_o[1][213] , \ootx_payload_o[1][214] , 
            \ootx_payload_o[1][215] , \ootx_payload_o[1][216] , \ootx_payload_o[1][217] , 
            \ootx_payload_o[1][218] , \ootx_payload_o[1][219] , \ootx_payload_o[1][220] , 
            \ootx_payload_o[1][221] , \ootx_payload_o[1][222] , \ootx_payload_o[1][223] , 
            \ootx_payload_o[1][224] , \ootx_payload_o[1][225] , \ootx_payload_o[1][226] , 
            \ootx_payload_o[1][227] , \ootx_payload_o[1][228] , \ootx_payload_o[1][229] , 
            \ootx_payload_o[1][230] , \ootx_payload_o[1][231] , \ootx_payload_o[1][232] , 
            \ootx_payload_o[1][233] , \ootx_payload_o[1][234] , \ootx_payload_o[1][235] , 
            \ootx_payload_o[1][236] , \ootx_payload_o[1][237] , \ootx_payload_o[1][238] , 
            \ootx_payload_o[1][239] , \ootx_payload_o[1][240] , \ootx_payload_o[1][241] , 
            \ootx_payload_o[1][242] , \ootx_payload_o[1][243] , \ootx_payload_o[1][244] , 
            \ootx_payload_o[1][245] , \ootx_payload_o[1][246] , \ootx_payload_o[1][247] , 
            \ootx_payload_o[1][248] , \ootx_payload_o[1][249] , \ootx_payload_o[1][250] , 
            \ootx_payload_o[1][251] , \ootx_payload_o[1][252] , \ootx_payload_o[1][253] , 
            \ootx_payload_o[1][254] , \ootx_payload_o[1][255] , \ootx_payload_o[1][256] , 
            \ootx_payload_o[1][257] , \ootx_payload_o[1][258] , \ootx_payload_o[1][259] , 
            \ootx_payload_o[1][260] , \ootx_payload_o[1][261] , \ootx_payload_o[1][262] , 
            \ootx_payload_o[1][263] , n860, n1264, ootx_payloads_1_215, 
            n586, n1401, ootx_payloads_1_214, n1359, ootx_payloads_1_213, 
            ootx_payloads_1_212, ootx_payloads_1_211, n584, n1402, n582, 
            n1403, ootx_payloads_1_210, n858, n1265, ootx_payloads_1_209, 
            n580, n1404, ootx_payloads_1_208, n578, n1405, n972, 
            n576, n1406, ootx_payloads_1_207, ootx_payloads_1_206, ootx_payloads_1_205, 
            ootx_payloads_1_204, ootx_payloads_1_203, n856, n1266, ootx_payloads_1_202, 
            n574, n1407, n970, n968, n572, n1408, ootx_payloads_1_201, 
            n854, n1267, n570, n1409, n740, n1324, ootx_payloads_1_200, 
            ootx_payloads_1_199, n738, n1325, n568, n1410, ootx_payloads_1_198, 
            n852, n1268, ootx_payloads_1_197, n566, n1411, ootx_payloads_1_196, 
            ootx_payloads_1_195, ootx_payloads_1_194, ootx_payloads_1_193, 
            ootx_payloads_1_192, n564, n1412, n850, n1269, n1360, 
            n562, n1413, n708, n1340, n560, n1414, n964, n9513, 
            ootx_payloads_N_1698, n558, n1415, ootx_payloads_1_191, 
            ootx_payloads_1_190, ootx_payloads_1_189, ootx_payloads_1_188, 
            ootx_payloads_1_187, n848, n1270, ootx_payloads_1_186, n556, 
            n1416, ootx_payloads_1_185, ootx_payloads_1_184, n554, n1417, 
            ootx_payloads_1_183, n768, n1310, n846, n1271, ootx_payloads_1_182, 
            n540, n542, n544, n546, n548, ootx_payloads_1_181, n550, 
            n552, n1370, n736, n686, n690, ootx_payloads_1_180, 
            n762, n692, ootx_payloads_1_179, n1313, n696, n698, 
            ootx_payloads_1_178, n700, n702, ootx_payloads_1_177, n936, 
            n1226, ootx_payloads_1_176, n704, ootx_payloads_1_175, ootx_payloads_1_174, 
            n706, ootx_payloads_1_173, ootx_payloads_1_172, ootx_payloads_1_171, 
            ootx_payloads_1_170, ootx_payloads_1_169, ootx_payloads_1_168, 
            ootx_payloads_1_167, ootx_payloads_1_166, ootx_payloads_1_165, 
            n962, ootx_payloads_1_164, ootx_payloads_1_163, ootx_payloads_1_162, 
            n646, n1371, ootx_payloads_1_161, ootx_payloads_1_160, n720, 
            ootx_payloads_1_159, n760, ootx_payloads_1_158, n1314, n642, 
            n644, ootx_payloads_1_157, ootx_payloads_1_156, ootx_payloads_1_155, 
            ootx_payloads_1_154, ootx_payloads_1_153, ootx_payloads_1_152, 
            ootx_payloads_1_151, ootx_payloads_1_150, ootx_payloads_1_149, 
            ootx_payloads_1_148, ootx_payloads_1_147, n960, ootx_payloads_1_146, 
            n770, n772, ootx_payloads_1_145, n774, n718, ootx_payloads_1_144, 
            ootx_payloads_1_143, n1361, n682, n684, ootx_payloads_1_142, 
            n688, ootx_payloads_1_141, ootx_payloads_1_140, n694, ootx_payloads_1_139, 
            ootx_payloads_1_138, ootx_payloads_1_137, ootx_payloads_1_136, 
            ootx_payloads_1_135, n734, n776, ootx_payloads_1_134, ootx_payloads_1_133, 
            ootx_payloads_1_132, ootx_payloads_1_131, n538, n756, n758, 
            ootx_payloads_1_130, ootx_payloads_1_129, n728, ootx_payloads_1_128, 
            ootx_payloads_1_127, n714, n730, n732, ootx_payloads_1_126, 
            ootx_payloads_1_125, ootx_payloads_1_124, ootx_payloads_1_123, 
            ootx_payloads_1_122, n716, ootx_payloads_1_121, ootx_payloads_1_120, 
            ootx_payloads_1_119, ootx_payloads_1_118, ootx_payloads_1_117, 
            ootx_payloads_1_116, ootx_payloads_1_115, n1315, ootx_payloads_1_114, 
            n722, ootx_payloads_1_113, ootx_payloads_1_112, ootx_payloads_1_111, 
            n1333, ootx_payloads_1_110, n726, ootx_payloads_1_109, ootx_payloads_1_108, 
            ootx_payloads_1_107, n1418, ootx_payloads_1_106, ootx_payloads_1_105, 
            ootx_payloads_1_104, ootx_payloads_1_103, ootx_payloads_1_102, 
            ootx_payloads_1_101, n1216, n844, n1272, n1217, ootx_payloads_1_100, 
            n1218, ootx_payloads_1_99, n1219, n842, n1273, n1419, 
            n1220, ootx_payloads_1_98, ootx_payloads_1_97, ootx_payloads_1_96, 
            n1221, ootx_payloads_1_95, ootx_payloads_1_94, ootx_payloads_1_93, 
            n1222, ootx_payloads_1_92, n1341, ootx_payloads_1_91, n1223, 
            ootx_payloads_1_90, n1224, ootx_payloads_1_89, ootx_payloads_1_88, 
            ootx_payloads_1_87, ootx_payloads_1_86, n840, n1274, ootx_payloads_1_85, 
            ootx_payloads_1_84, ootx_payloads_1_83, n1420, n1227, ootx_payloads_1_82, 
            n1228, n838, n1275, ootx_payloads_1_81, n934, n1229, 
            ootx_payloads_1_80, ootx_payloads_1_79, ootx_payloads_1_78, 
            ootx_payloads_1_77, ootx_payloads_1_76, ootx_payloads_1_75, 
            n1342, n1421, ootx_payloads_1_74, n836, n1276, ootx_payloads_1_73, 
            ootx_payloads_1_72, n1422, n1423, n834, n1277, ootx_payloads_1_71, 
            ootx_payloads_1_70, n1424, ootx_payloads_1_69, ootx_payloads_1_68, 
            ootx_payloads_1_67, ootx_payloads_1_66, ootx_payloads_1_65, 
            ootx_payloads_1_64, n1343, n1425, ootx_payloads_1_63, n832, 
            n1278, ootx_payloads_1_62, ootx_payloads_1_61, n536, n1426, 
            n1316, ootx_payloads_1_60, n1334, ootx_payloads_1_59, ootx_payloads_1_58, 
            ootx_payloads_1_57, n534, n1427, ootx_payloads_1_56, n830, 
            n1279, n1362, ootx_payloads_1_55, ootx_payloads_1_54, ootx_payloads_1_53, 
            n1344, n532, n1428, ootx_payloads_1_52, n828, n1280, 
            n530, n1429, n956, n1345, ootx_payloads_1_51, ootx_payloads_1_50, 
            ootx_payloads_1_49, n954, n826, n1281, ootx_payloads_1_48, 
            n528, n1430, ootx_payloads_1_47, n526, n1431, ootx_payloads_1_46, 
            ootx_payloads_1_45, n1346, n824, n1282, ootx_payloads_1_44, 
            n952, ootx_payloads_1_43, n524, n1432, \ootx_payloads_N_1730[12] , 
            ootx_payloads_1_42, ootx_payloads_1_41, ootx_payloads_1_40, 
            ootx_payloads_1_39, ootx_payloads_1_38, ootx_payloads_1_37, 
            n522, n1433, n822, n1283, n1347, n950, \ootx_payloads_N_1730[11] , 
            ootx_payloads_1_36, ootx_payloads_1_35, n1326, ootx_payloads_1_34, 
            ootx_payloads_1_33, n1348, n6334, ootx_payloads_1_32, ootx_payloads_1_31, 
            n51, n52, ootx_payloads_1_30, n948, \ootx_payloads_N_1730[10] , 
            ootx_payloads_1_29, ootx_payloads_1_28, n2679, n2680, n6335, 
            n1349, ootx_payloads_1_27, n1317, n932, ootx_payloads_1_26, 
            n6336, n946, ootx_payloads_1_25, ootx_payloads_1_24, ootx_payloads_1_23, 
            \ootx_payloads_N_1730[9] , n1363, ootx_payloads_1_22, n49, 
            n50, n9771, n820, n1284, ootx_payloads_1_21, n6337, 
            ootx_payloads_1_20, n1350, ootx_payloads_1_19, ootx_payloads_1_18, 
            ootx_payloads_1_17, n944, n6338, ootx_payloads_1_16, n1351, 
            \ootx_payloads_N_1730[8] , n47, n48, n818, n1285, ootx_payloads_1_15, 
            ootx_payloads_1_14, ootx_payloads_1_13, ootx_payloads_1_12, 
            n942, n6339, ootx_payloads_1_11, n45, n46, ootx_payloads_1_10, 
            \ootx_payloads_N_1730[7] , n816, n1286, ootx_payloads_1_9, 
            n6340, ootx_payloads_1_8, crc32s_1_25, crc32s_1_30, crc32s_1_27, 
            crc32s_1_26, crc32s_1_31, crc32s_1_29, crc32s_1_28, crc32s_1_24, 
            crc32s_1_23, crc32s_1_22, crc32s_1_21, ootx_payloads_1_7, 
            crc32s_1_20, \ootx_payloads_N_1730[6] , n1364, ootx_payloads_1_6, 
            ootx_payloads_1_5, crc32s_1_19, crc32s_1_18, crc32s_1_17, 
            crc32s_1_16, crc32s_1_15, n6341, crc32s_1_14, crc32s_1_13, 
            crc32s_1_12, crc32s_1_11, crc32s_1_10, crc32s_1_9, crc32s_1_8, 
            crc32s_1_7, crc32s_1_6, crc32s_1_5, crc32s_1_4, crc32s_1_3, 
            crc32s_1_2, ootx_payloads_1_4, ootx_payloads_1_3, crc32s_1_0, 
            ootx_payloads_1_2, crc32s_1_1, \ootx_payloads_N_1730[5] , 
            ootx_payloads_1_1, n43, n6342, n44, n28, n814, n1287, 
            n41, n42, n1288, n1289, n1290, n1291, n1292, n1293, 
            n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
            n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
            n1327, n1328, n1329, n1330, n1331, n1335, n1336, n1337, 
            n1352, n1353, n1365, n1366, n1367, n1368, n1369, n1372, 
            n1373, n11612, n3112, n11611, n11610, n11609, n11608, 
            n11607, n11606, n11605, n11604, n22997, n11602, n23001, 
            n11600, n11599, n11598, n11597, n11596, n11595, n11594, 
            n11593, n11592, n11591, n11590, n11589, n11588, n11587, 
            n11586, n11585, n11584, n11583, n11582, n11581, n11580, 
            n11579, n11578, n11577, n11576, n11575, n11574, n11573, 
            n11572, n11571, n11570, n11569, n11568, n11567, n11566, 
            n11565, n11564, n11563, n11562, n11561, n11560, n11559, 
            n11558, n11557, n11556, n11555, n11554, n11553, n11552, 
            n11551, n11550, n11549, n11548, n11547, n11546, n11545, 
            n11544, n11543, n11542, n11541, n11540, n11539, n11538, 
            n11537, n11536, n11535, n11534, n11533, n11532, n11531, 
            n11530, n11529, n11528, n11527, n11526, n11525, n11524, 
            n11523, n11522, n11521, n11520, n11519, n11518, n11517, 
            n11516, n11515, n11514, n11513, n11512, n11511, n11510, 
            n11509, n11508, n11507, n11506, n11505, n11504, n39, 
            n40, n812, n37, n38, n6343, n810, n808, n17, n19468, 
            n806, n535, n792, n804, n533, led_c_0, n790, led_c_1, 
            led_c_2, led_c_3, led_c_4, led_c_5, led_c_6, n802, n800, 
            n531, n11503, n11502, n11501, n11500, n11499, n11498, 
            n11497, n11496, n11495, n11494, n11493, n11492, n11491, 
            n11490, n11489, n11488, n11487, n11486, n11485, n11484, 
            n11483, n11482, n11481, n11480, n11479, n11478, n11477, 
            n11476, n11475, n11474, n11473, n11472, n788, n11471, 
            n11470, n11469, n11468, n11467, n11466, n11465, n11464, 
            n11463, n11462, n11461, n11460, n11459, n11458, n11457, 
            n11456, n11455, n11454, n11453, n11452, n11451, n11450, 
            n11449, n11448, n11447, n11446, n11445, n11444, n11443, 
            n11442, n11441, n11440, n11439, n11438, n11437, n11436, 
            n11435, n11434, n11433, n11432, n11431, n11430, n11429, 
            n11428, n11427, n11426, n11425, n11424, n11423, n11422, 
            n11421, n11420, n11419, n11418, n11417, n11416, n11415, 
            n11414, n11413, n11412, n11411, n11410, n11409, n11408, 
            n11407, n11406, n11405, n11404, n11403, n11402, n11401, 
            n11400, n11399, n11398, n11397, n11396, n11395, n11394, 
            n11393, n11392, n11391, n11390, n11389, n11388, n11387, 
            n11386, n11385, n11384, n11383, n11382, n11381, n11380, 
            n11379, n11378, n11377, n11376, n11375, n11374, n11373, 
            n11372, n11371, n11370, n11369, n11368, n11367, n11366, 
            n11365, n11364, n11363, n11362, n11361, n11360, n11359, 
            n11358, n11357, n11356, n11355, n11354, n11353, n11352, 
            n11351, n11350, n11349, n11348, n11347, n11346, n11345, 
            n11344, n11343, n11342, n11341, n11340, n11339, n11338, 
            n11337, n11336, n11335, n11334, n11333, n11332, n11331, 
            n11330, n11329, n11328, n11327, n11326, n11325, n11324, 
            n11323, n11322, n11321, n11320, n11319, n11318, n11317, 
            n11316, n11315, n11314, n11313, n11312, n11311, n11310, 
            n11309, n11308, n11307, n11306, n11305, n11304, n11303, 
            n11302, n11301, n11300, n11299, n11298, n11297, n11296, 
            n11295, n11294, n11293, n11292, n11291, n11290, n11289, 
            n11288, n11287, n11286, n11285, ootx_payloads_1_0, n6344, 
            n798, n529, n796, n6345, n786, n794, n527, n6346, 
            n784, n525, n782, n523, n780, n778, n521, n1032, 
            \ootx_payloads_N_1730[0] , n930, n940, sync, n1022, n1012, 
            n1014, n1002, n1016, n1018, n1020, n1024, n1026, n1028, 
            n1030, n11016, \ootx_payload_o[0][0] , n67, n65, n63, 
            \ootx_states[1][0] , n25, n61, n59, n57, n55, n53, 
            n68, n66, n64, n62, n60, n58, n56, n54, n20_adj_33, 
            led_c_7);
    output \lighthouse[0] ;
    output [31:0]n6333;
    output [31:0]counter_from_last_rise;
    input GND_net;
    output \ootx_payload_o[1][0] ;
    input clock_c;
    output n1;
    output n1_adj_1;
    output n1000;
    output data;
    output n1194;
    output \ootx_payloads_N_1730[1] ;
    output [30:0]n2851;
    output bit_counters_0_7;
    output bit_counters_1_7;
    output bit_counters_0_8;
    output bit_counters_1_8;
    output bit_counters_0_9;
    output bit_counters_1_9;
    output \ootx_payloads_N_1730[2] ;
    output n24018;
    output \ootx_payloads_N_1699[4] ;
    output n13221;
    input reset_c;
    output new_data;
    output [1:0]ootx_payloads_N_1744;
    output bit_counters_0_10;
    output bit_counters_1_10;
    output \ootx_payloads_N_1730[3] ;
    output [30:0]n337;
    output n998;
    output n1195;
    output n996;
    output n1196;
    output n994;
    output n1197;
    input VCC_net;
    output n992;
    output n1198;
    output n766;
    output n1311;
    output n13;
    output n990;
    output n1199;
    output n988;
    output n1200;
    output n1_adj_2;
    output n9797;
    input n23974;
    input n8;
    output bit_counters_0_19;
    output bit_counters_1_19;
    input n23003;
    output data_counters_0_0;
    input n23005;
    output data_counters_0_1;
    input n23007;
    output data_counters_0_2;
    input n23009;
    output data_counters_0_3;
    input n23011;
    output data_counters_0_4;
    input n23013;
    output data_counters_0_5;
    input n23015;
    output data_counters_0_6;
    input n23017;
    output data_counters_0_7;
    input n23019;
    output data_counters_0_8;
    input n23021;
    output data_counters_0_9;
    input n23023;
    output data_counters_0_10;
    output n1_adj_3;
    input n23025;
    output data_counters_0_11;
    input n23027;
    output data_counters_0_12;
    input n23029;
    output data_counters_0_13;
    input n23031;
    output data_counters_0_14;
    input n23033;
    output data_counters_0_15;
    input n23035;
    output data_counters_0_16;
    input n23037;
    output data_counters_0_17;
    input n23039;
    output data_counters_0_18;
    input n23041;
    output data_counters_0_19;
    input n23043;
    output data_counters_0_20;
    input n23045;
    output data_counters_0_21;
    input n23047;
    output data_counters_0_22;
    input n23049;
    output data_counters_0_23;
    input n23051;
    output data_counters_0_24;
    input n23053;
    output data_counters_0_25;
    input n23055;
    output data_counters_0_26;
    input n23057;
    output data_counters_0_27;
    input n23059;
    output data_counters_0_28;
    input n23061;
    output data_counters_0_29;
    input n23063;
    output data_counters_0_30;
    input n23065;
    output data_counters_1_0;
    input n23067;
    output data_counters_1_1;
    input n23069;
    output data_counters_1_2;
    input n23071;
    output data_counters_1_3;
    input n23073;
    output data_counters_1_4;
    input n23075;
    output data_counters_1_5;
    input n23077;
    output data_counters_1_6;
    input n23079;
    output data_counters_1_7;
    input n23081;
    output data_counters_1_8;
    input n23083;
    output data_counters_1_9;
    input n23085;
    output data_counters_1_10;
    input n23087;
    output data_counters_1_11;
    input n23089;
    output data_counters_1_12;
    input n23091;
    output data_counters_1_13;
    input n23093;
    output data_counters_1_14;
    input n23095;
    output data_counters_1_15;
    input n23097;
    output data_counters_1_16;
    input n23099;
    output data_counters_1_17;
    input n23101;
    output data_counters_1_18;
    input n23103;
    output data_counters_1_19;
    input n23105;
    output data_counters_1_20;
    input n23107;
    output data_counters_1_21;
    input n23109;
    output data_counters_1_22;
    input n23111;
    output data_counters_1_23;
    input n23113;
    output data_counters_1_24;
    input n23115;
    output data_counters_1_25;
    input n23117;
    output data_counters_1_26;
    input n23119;
    output data_counters_1_27;
    input n23121;
    output data_counters_1_28;
    input n23123;
    output data_counters_1_29;
    input n23125;
    output data_counters_1_30;
    input n23475;
    output bit_counters_0_0;
    input n23477;
    output bit_counters_0_1;
    input n23479;
    output bit_counters_0_2;
    input n23481;
    output bit_counters_0_3;
    input n23483;
    output bit_counters_0_4;
    input n23485;
    output bit_counters_0_5;
    input n23487;
    output bit_counters_0_6;
    input n23489;
    input n23491;
    input n23493;
    input n23495;
    input n23497;
    output bit_counters_0_11;
    input n23499;
    output bit_counters_0_12;
    input n23501;
    output bit_counters_0_13;
    input n23503;
    output bit_counters_0_14;
    input n23505;
    output bit_counters_0_15;
    input n23507;
    output bit_counters_0_16;
    input n23509;
    output bit_counters_0_17;
    input n23469;
    output bit_counters_0_18;
    input n23463;
    input n23457;
    output bit_counters_0_20;
    input n23451;
    output bit_counters_0_21;
    input n23445;
    output bit_counters_0_22;
    input n23439;
    output bit_counters_0_23;
    input n23433;
    output bit_counters_0_24;
    input n23427;
    output bit_counters_0_25;
    input n23421;
    output bit_counters_0_26;
    input n23415;
    output bit_counters_0_27;
    input n23409;
    output bit_counters_0_28;
    input n23399;
    output bit_counters_0_29;
    input n23389;
    output bit_counters_0_30;
    input n23511;
    output bit_counters_1_0;
    input n23513;
    output bit_counters_1_1;
    input n23515;
    output bit_counters_1_2;
    input n23517;
    output bit_counters_1_3;
    input n23519;
    output bit_counters_1_4;
    input n23521;
    output bit_counters_1_5;
    input n23523;
    output bit_counters_1_6;
    input n23525;
    input n23527;
    input n23529;
    input n23531;
    input n23533;
    output bit_counters_1_11;
    input n23535;
    output bit_counters_1_12;
    input n23537;
    output bit_counters_1_13;
    input n23539;
    output bit_counters_1_14;
    input n23541;
    output bit_counters_1_15;
    input n23543;
    output bit_counters_1_16;
    input n23545;
    output bit_counters_1_17;
    input n23471;
    output bit_counters_1_18;
    input n23465;
    input n23459;
    output bit_counters_1_20;
    input n23453;
    output bit_counters_1_21;
    input n23447;
    output bit_counters_1_22;
    input n23441;
    output bit_counters_1_23;
    input n23435;
    output bit_counters_1_24;
    input n23429;
    output bit_counters_1_25;
    input n23423;
    output bit_counters_1_26;
    input n23417;
    output bit_counters_1_27;
    output n986;
    output n1201;
    output n35;
    input n23411;
    output bit_counters_1_28;
    input n23401;
    output bit_counters_1_29;
    input n23391;
    output bit_counters_1_30;
    input n23697;
    input n23639;
    output payload_lengths_0_0;
    input n23641;
    output payload_lengths_1_0;
    input n8_adj_4;
    input n8_adj_5;
    input n8_adj_6;
    output n2282;
    input n8_adj_7;
    output n984;
    output n1202;
    input n8_adj_8;
    output \counter_from_last_rise[6] ;
    input n8_adj_9;
    output \counter_from_last_rise[7] ;
    input n8_adj_10;
    output \counter_from_last_rise[8] ;
    input n8_adj_11;
    output \counter_from_last_rise[9] ;
    input n8_adj_12;
    output \counter_from_last_rise[10] ;
    input n8_adj_13;
    output \counter_from_last_rise[11] ;
    input n8_adj_14;
    output \counter_from_last_rise[12] ;
    input n8_adj_15;
    input n8_adj_16;
    input n8_adj_17;
    input n8_adj_18;
    input n8_adj_19;
    input n8_adj_20;
    input n8_adj_21;
    output \counter_from_last_rise[19] ;
    input n8_adj_22;
    output \counter_from_last_rise[20] ;
    input n8_adj_23;
    output \counter_from_last_rise[21] ;
    input n8_adj_24;
    output \counter_from_last_rise[22] ;
    input n8_adj_25;
    output \counter_from_last_rise[23] ;
    input n8_adj_26;
    output \counter_from_last_rise[24] ;
    input n8_adj_27;
    output \counter_from_last_rise[25] ;
    input n8_adj_28;
    output \counter_from_last_rise[26] ;
    input n8_adj_29;
    output \counter_from_last_rise[27] ;
    input n8_adj_30;
    output \counter_from_last_rise[28] ;
    input n8_adj_31;
    output \counter_from_last_rise[29] ;
    input n23407;
    output \counter_from_last_rise[30] ;
    input n23397;
    output \counter_from_last_rise[31] ;
    input n12201;
    output \ootx_payload_o[0][263] ;
    input n12200;
    output \ootx_payload_o[0][262] ;
    input n12199;
    output \ootx_payload_o[0][261] ;
    input n12198;
    output \ootx_payload_o[0][260] ;
    input n12197;
    output \ootx_payload_o[0][259] ;
    input n12196;
    output \ootx_payload_o[0][258] ;
    input n12195;
    output \ootx_payload_o[0][257] ;
    input n12194;
    output \ootx_payload_o[0][256] ;
    input n12193;
    output \ootx_payload_o[0][255] ;
    input n12192;
    output \ootx_payload_o[0][254] ;
    input n12191;
    output \ootx_payload_o[0][253] ;
    input n12190;
    output \ootx_payload_o[0][252] ;
    input n12189;
    output \ootx_payload_o[0][251] ;
    input n12188;
    output \ootx_payload_o[0][250] ;
    input n12187;
    output \ootx_payload_o[0][249] ;
    input n12186;
    output \ootx_payload_o[0][248] ;
    input n12185;
    output \ootx_payload_o[0][247] ;
    input n12184;
    output \ootx_payload_o[0][246] ;
    input n12183;
    output \ootx_payload_o[0][245] ;
    input n12182;
    output \ootx_payload_o[0][244] ;
    input n12181;
    output \ootx_payload_o[0][243] ;
    input n12180;
    output \ootx_payload_o[0][242] ;
    input n12179;
    output \ootx_payload_o[0][241] ;
    input n12178;
    output \ootx_payload_o[0][240] ;
    input n12177;
    output \ootx_payload_o[0][239] ;
    input n12176;
    output \ootx_payload_o[0][238] ;
    input n12175;
    output \ootx_payload_o[0][237] ;
    input n12174;
    output \ootx_payload_o[0][236] ;
    input n12173;
    output \ootx_payload_o[0][235] ;
    input n12172;
    output \ootx_payload_o[0][234] ;
    input n12171;
    output \ootx_payload_o[0][233] ;
    input n12170;
    output \ootx_payload_o[0][232] ;
    input n12169;
    output \ootx_payload_o[0][231] ;
    input n12168;
    output \ootx_payload_o[0][230] ;
    input n12167;
    output \ootx_payload_o[0][229] ;
    input n12166;
    output \ootx_payload_o[0][228] ;
    input n12165;
    output \ootx_payload_o[0][227] ;
    input n12164;
    output \ootx_payload_o[0][226] ;
    input n12163;
    output \ootx_payload_o[0][225] ;
    input n12162;
    output \ootx_payload_o[0][224] ;
    input n12161;
    output \ootx_payload_o[0][223] ;
    input n12160;
    output \ootx_payload_o[0][222] ;
    input n12159;
    output \ootx_payload_o[0][221] ;
    input n12158;
    output \ootx_payload_o[0][220] ;
    input n12157;
    output \ootx_payload_o[0][219] ;
    input n12156;
    output \ootx_payload_o[0][218] ;
    input n12155;
    output \ootx_payload_o[0][217] ;
    input n12154;
    output \ootx_payload_o[0][216] ;
    input n12153;
    output \ootx_payload_o[0][215] ;
    input n12152;
    output \ootx_payload_o[0][214] ;
    input n12151;
    output \ootx_payload_o[0][213] ;
    input n12150;
    output \ootx_payload_o[0][212] ;
    input n12149;
    output \ootx_payload_o[0][211] ;
    input n12148;
    output \ootx_payload_o[0][210] ;
    input n12147;
    output \ootx_payload_o[0][209] ;
    input n12146;
    output \ootx_payload_o[0][208] ;
    input n12145;
    output \ootx_payload_o[0][207] ;
    input n12144;
    output \ootx_payload_o[0][206] ;
    input n12143;
    output \ootx_payload_o[0][205] ;
    input n12142;
    output \ootx_payload_o[0][204] ;
    input n12141;
    output \ootx_payload_o[0][203] ;
    input n12140;
    output \ootx_payload_o[0][202] ;
    input n12139;
    output \ootx_payload_o[0][201] ;
    input n12138;
    output \ootx_payload_o[0][200] ;
    input n12137;
    output \ootx_payload_o[0][199] ;
    input n12136;
    output \ootx_payload_o[0][198] ;
    input n12135;
    output \ootx_payload_o[0][197] ;
    input n12134;
    output \ootx_payload_o[0][196] ;
    input n12133;
    output \ootx_payload_o[0][195] ;
    input n12132;
    output \ootx_payload_o[0][194] ;
    input n12131;
    output \ootx_payload_o[0][193] ;
    input n12130;
    output \ootx_payload_o[0][192] ;
    input n12129;
    output \ootx_payload_o[0][191] ;
    input n12128;
    output \ootx_payload_o[0][190] ;
    input n12127;
    output \ootx_payload_o[0][189] ;
    input n12126;
    output \ootx_payload_o[0][188] ;
    input n12125;
    output \ootx_payload_o[0][187] ;
    input n12124;
    output \ootx_payload_o[0][186] ;
    input n12123;
    output \ootx_payload_o[0][185] ;
    input n12122;
    output \ootx_payload_o[0][184] ;
    input n12121;
    output \ootx_payload_o[0][183] ;
    input n12120;
    output \ootx_payload_o[0][182] ;
    input n12119;
    output \ootx_payload_o[0][181] ;
    input n12118;
    output \ootx_payload_o[0][180] ;
    input n12117;
    output \ootx_payload_o[0][179] ;
    input n12116;
    output \ootx_payload_o[0][178] ;
    input n12115;
    output \ootx_payload_o[0][177] ;
    input n12114;
    output \ootx_payload_o[0][176] ;
    input n12113;
    output \ootx_payload_o[0][175] ;
    input n12112;
    output \ootx_payload_o[0][174] ;
    input n12111;
    output \ootx_payload_o[0][173] ;
    input n12110;
    output \ootx_payload_o[0][172] ;
    input n12109;
    output \ootx_payload_o[0][171] ;
    input n12108;
    output \ootx_payload_o[0][170] ;
    input n12107;
    output \ootx_payload_o[0][169] ;
    input n12106;
    output \ootx_payload_o[0][168] ;
    input n12105;
    output \ootx_payload_o[0][167] ;
    input n12104;
    output \ootx_payload_o[0][166] ;
    input n12103;
    output \ootx_payload_o[0][165] ;
    input n12102;
    output \ootx_payload_o[0][164] ;
    input n12101;
    output \ootx_payload_o[0][163] ;
    input n12100;
    output \ootx_payload_o[0][162] ;
    input n12099;
    output \ootx_payload_o[0][161] ;
    input n12098;
    output \ootx_payload_o[0][160] ;
    input n12097;
    output \ootx_payload_o[0][159] ;
    input n12096;
    output \ootx_payload_o[0][158] ;
    input n12095;
    output \ootx_payload_o[0][157] ;
    input n12094;
    output \ootx_payload_o[0][156] ;
    input n12093;
    output \ootx_payload_o[0][155] ;
    input n12092;
    output \ootx_payload_o[0][154] ;
    input n12091;
    output \ootx_payload_o[0][153] ;
    input n12090;
    output \ootx_payload_o[0][152] ;
    input n12089;
    output \ootx_payload_o[0][151] ;
    input n12088;
    output \ootx_payload_o[0][150] ;
    input n12087;
    output \ootx_payload_o[0][149] ;
    input n12086;
    output \ootx_payload_o[0][148] ;
    input n12085;
    output \ootx_payload_o[0][147] ;
    input n12084;
    output \ootx_payload_o[0][146] ;
    input n12083;
    output \ootx_payload_o[0][145] ;
    input n12082;
    output \ootx_payload_o[0][144] ;
    input n12081;
    output \ootx_payload_o[0][143] ;
    input n12080;
    output \ootx_payload_o[0][142] ;
    input n12079;
    output \ootx_payload_o[0][141] ;
    input n12078;
    output \ootx_payload_o[0][140] ;
    input n12077;
    output \ootx_payload_o[0][139] ;
    input n12076;
    output \ootx_payload_o[0][138] ;
    input n12075;
    output \ootx_payload_o[0][137] ;
    input n12074;
    output \ootx_payload_o[0][136] ;
    input n12073;
    output \ootx_payload_o[0][135] ;
    input n12072;
    output \ootx_payload_o[0][134] ;
    input n12071;
    output \ootx_payload_o[0][133] ;
    input n12070;
    output \ootx_payload_o[0][132] ;
    input n12069;
    output \ootx_payload_o[0][131] ;
    input n12068;
    output \ootx_payload_o[0][130] ;
    input n12067;
    output \ootx_payload_o[0][129] ;
    input n12066;
    output \ootx_payload_o[0][128] ;
    input n12065;
    output \ootx_payload_o[0][127] ;
    input n12064;
    output \ootx_payload_o[0][126] ;
    input n12063;
    output \ootx_payload_o[0][125] ;
    input n12062;
    output \ootx_payload_o[0][124] ;
    input n12061;
    output \ootx_payload_o[0][123] ;
    input n12060;
    output \ootx_payload_o[0][122] ;
    input n12059;
    output \ootx_payload_o[0][121] ;
    input n12058;
    output \ootx_payload_o[0][120] ;
    input n12057;
    output \ootx_payload_o[0][119] ;
    input n12056;
    output \ootx_payload_o[0][118] ;
    input n12055;
    output \ootx_payload_o[0][117] ;
    input n12054;
    output \ootx_payload_o[0][116] ;
    input n12053;
    output \ootx_payload_o[0][115] ;
    input n12052;
    output \ootx_payload_o[0][114] ;
    input n12051;
    output \ootx_payload_o[0][113] ;
    input n12050;
    output \ootx_payload_o[0][112] ;
    input n12049;
    output \ootx_payload_o[0][111] ;
    input n12048;
    output \ootx_payload_o[0][110] ;
    input n12047;
    output \ootx_payload_o[0][109] ;
    input n12046;
    output \ootx_payload_o[0][108] ;
    input n12045;
    output \ootx_payload_o[0][107] ;
    input n12044;
    output \ootx_payload_o[0][106] ;
    input n12043;
    output \ootx_payload_o[0][105] ;
    input n12042;
    output \ootx_payload_o[0][104] ;
    input n12041;
    output \ootx_payload_o[0][103] ;
    input n12040;
    output \ootx_payload_o[0][102] ;
    input n12039;
    output \ootx_payload_o[0][101] ;
    input n12038;
    output \ootx_payload_o[0][100] ;
    input n12037;
    output \ootx_payload_o[0][99] ;
    input n12036;
    output \ootx_payload_o[0][98] ;
    input n12035;
    output \ootx_payload_o[0][97] ;
    input n12034;
    output \ootx_payload_o[0][96] ;
    input n12033;
    output \ootx_payload_o[0][95] ;
    input n12032;
    output \ootx_payload_o[0][94] ;
    input n12031;
    output \ootx_payload_o[0][93] ;
    input n12030;
    output \ootx_payload_o[0][92] ;
    input n12029;
    output \ootx_payload_o[0][91] ;
    input n12028;
    output \ootx_payload_o[0][90] ;
    input n12027;
    output \ootx_payload_o[0][89] ;
    input n12026;
    output \ootx_payload_o[0][88] ;
    input n12025;
    output \ootx_payload_o[0][87] ;
    input n12024;
    output \ootx_payload_o[0][86] ;
    input n12023;
    output \ootx_payload_o[0][85] ;
    input n12022;
    output \ootx_payload_o[0][84] ;
    input n12021;
    output \ootx_payload_o[0][83] ;
    input n12020;
    output \ootx_payload_o[0][82] ;
    input n12019;
    output \ootx_payload_o[0][81] ;
    input n12018;
    output \ootx_payload_o[0][80] ;
    input n12017;
    output \ootx_payload_o[0][79] ;
    input n12016;
    output \ootx_payload_o[0][78] ;
    input n12015;
    output \ootx_payload_o[0][77] ;
    input n12014;
    output \ootx_payload_o[0][76] ;
    input n12013;
    output \ootx_payload_o[0][75] ;
    input n12012;
    output \ootx_payload_o[0][74] ;
    input n12011;
    output \ootx_payload_o[0][73] ;
    input n12010;
    output \ootx_payload_o[0][72] ;
    input n12009;
    output \ootx_payload_o[0][71] ;
    input n12008;
    output \ootx_payload_o[0][70] ;
    input n12007;
    output \ootx_payload_o[0][69] ;
    input n12006;
    output \ootx_payload_o[0][68] ;
    input n12005;
    output \ootx_payload_o[0][67] ;
    input n12004;
    output \ootx_payload_o[0][66] ;
    input n12003;
    output \ootx_payload_o[0][65] ;
    input n12002;
    output \ootx_payload_o[0][64] ;
    input n12001;
    output \ootx_payload_o[0][63] ;
    input n12000;
    output \ootx_payload_o[0][62] ;
    input n11999;
    output \ootx_payload_o[0][61] ;
    input n11998;
    output \ootx_payload_o[0][60] ;
    input n11997;
    output \ootx_payload_o[0][59] ;
    input n11996;
    output \ootx_payload_o[0][58] ;
    input n11995;
    output \ootx_payload_o[0][57] ;
    input n11994;
    output \ootx_payload_o[0][56] ;
    input n11993;
    output \ootx_payload_o[0][55] ;
    input n11992;
    output \ootx_payload_o[0][54] ;
    input n11991;
    output \ootx_payload_o[0][53] ;
    input n11990;
    output \ootx_payload_o[0][52] ;
    output n938;
    output n1225;
    input n11989;
    output \ootx_payload_o[0][51] ;
    input n11988;
    output \ootx_payload_o[0][50] ;
    input n11987;
    output \ootx_payload_o[0][49] ;
    input n11986;
    output \ootx_payload_o[0][48] ;
    input n11985;
    output \ootx_payload_o[0][47] ;
    input n11984;
    output \ootx_payload_o[0][46] ;
    input n11983;
    output \ootx_payload_o[0][45] ;
    output n958;
    output n1215;
    input n11982;
    output \ootx_payload_o[0][44] ;
    input n30;
    input n11981;
    output \ootx_payload_o[0][43] ;
    input n11980;
    output \ootx_payload_o[0][42] ;
    input n11979;
    output \ootx_payload_o[0][41] ;
    input n11978;
    output \ootx_payload_o[0][40] ;
    input n11977;
    output \ootx_payload_o[0][39] ;
    output n982;
    output n1203;
    input n11976;
    output \ootx_payload_o[0][38] ;
    input n11975;
    output \ootx_payload_o[0][37] ;
    input n11974;
    output \ootx_payload_o[0][36] ;
    input n11973;
    output \ootx_payload_o[0][35] ;
    output sensor_state;
    input n11972;
    output \ootx_payload_o[0][34] ;
    input n11971;
    output \ootx_payload_o[0][33] ;
    input n11970;
    output \ootx_payload_o[0][32] ;
    input n11969;
    output \ootx_payload_o[0][31] ;
    input n11968;
    output \ootx_payload_o[0][30] ;
    input n11967;
    output \ootx_payload_o[0][29] ;
    input n11966;
    output \ootx_payload_o[0][28] ;
    input n11965;
    output \ootx_payload_o[0][27] ;
    input n11964;
    output \ootx_payload_o[0][26] ;
    input n11963;
    output \ootx_payload_o[0][25] ;
    input n11962;
    output \ootx_payload_o[0][24] ;
    input n11961;
    output \ootx_payload_o[0][23] ;
    input n11960;
    output \ootx_payload_o[0][22] ;
    input n11959;
    output \ootx_payload_o[0][21] ;
    output n680;
    output n1354;
    output n712;
    output n1338;
    output \ootx_payloads_N_1699[5] ;
    output \ootx_payloads_N_1699[3] ;
    output \ootx_payloads_N_1699[15] ;
    output [1:0]n34;
    input n11958;
    output \ootx_payload_o[0][20] ;
    input n11957;
    output \ootx_payload_o[0][19] ;
    input n11956;
    output \ootx_payload_o[0][18] ;
    input n11955;
    output \ootx_payload_o[0][17] ;
    input n11954;
    output \ootx_payload_o[0][16] ;
    input n11953;
    output \ootx_payload_o[0][15] ;
    input n11952;
    output \ootx_payload_o[0][14] ;
    input n11951;
    output \ootx_payload_o[0][13] ;
    input n11950;
    output \ootx_payload_o[0][12] ;
    input n11949;
    output \ootx_payload_o[0][11] ;
    input n11948;
    output \ootx_payload_o[0][10] ;
    input n11947;
    output \ootx_payload_o[0][9] ;
    input n11946;
    output \ootx_payload_o[0][8] ;
    input n11945;
    output \ootx_payload_o[0][7] ;
    input n11944;
    output \ootx_payload_o[0][6] ;
    input n11943;
    output \ootx_payload_o[0][5] ;
    input n11942;
    output \ootx_payload_o[0][4] ;
    input n11941;
    output \ootx_payload_o[0][3] ;
    input n11940;
    output \ootx_payload_o[0][2] ;
    input n11939;
    output \ootx_payload_o[0][1] ;
    output [31:0]\ootx_crc32_o[1] ;
    output [31:0]\ootx_crc32_o[0] ;
    output n1170;
    output n1171;
    output n1172;
    output n1173;
    output n1174;
    output n1175;
    output n1176;
    output n1177;
    output n1178;
    output n1179;
    output n1180;
    output n1181;
    output n1182;
    output n1183;
    output n1184;
    output n1185;
    output n1186;
    output n1187;
    output n1188;
    output n1189;
    output n1190;
    output n1191;
    output n1192;
    output n1193;
    output n640;
    output n1374;
    output n724;
    output n928;
    output n1230;
    output n1204;
    output n1205;
    output n1206;
    output n1207;
    output n1208;
    output n1209;
    output n1210;
    output n1332;
    output n1211;
    output n1212;
    output n1213;
    output \ootx_payloads_N_1699[6] ;
    output \ootx_payloads_N_1699[7] ;
    output \ootx_payloads_N_1699[8] ;
    output n1010;
    output n1214;
    output n754;
    output n764;
    output n672;
    output [1:0]\ootx_states[0] ;
    output n638;
    output n1375;
    output ootx_payloads_1_263;
    output n926;
    output n1231;
    output n670;
    output n1312;
    output n20;
    output ootx_payloads_1_262;
    output n924;
    output n1232;
    output n636;
    output n1376;
    output n668;
    output n922;
    output n1233;
    output n634;
    output n1377;
    output n666;
    output n920;
    output n1234;
    output n632;
    output n1378;
    output n664;
    output n918;
    output n1235;
    output n662;
    output n916;
    output n1236;
    output n752;
    output n1318;
    output n660;
    output n914;
    output n1237;
    output n658;
    output n678;
    output n1355;
    output n912;
    output n1238;
    output n630;
    output n1379;
    output ootx_payloads_1_261;
    output ootx_payloads_1_260;
    output n656;
    output ootx_payloads_1_259;
    output n910;
    output n1239;
    output n654;
    output n1008;
    output n676;
    output n1356;
    output n908;
    output n1240;
    output ootx_payloads_1_258;
    output ootx_payloads_1_257;
    output ootx_payloads_1_256;
    output n628;
    output n1380;
    output ootx_payloads_1_255;
    output \ootx_payloads_N_1699[30] ;
    output n9200;
    output \ootx_payloads_N_1699[9] ;
    output \ootx_payloads_N_1699[13] ;
    output \ootx_payloads_N_1699[12] ;
    output \ootx_payloads_N_1699[11] ;
    output ootx_payloads_1_254;
    output ootx_payloads_1_253;
    output ootx_payloads_1_252;
    output ootx_payloads_1_251;
    output n652;
    output n906;
    output n1241;
    output ootx_payloads_1_250;
    output ootx_payloads_1_249;
    output \ootx_payloads_N_1699[10] ;
    output \ootx_payloads_N_1699[14] ;
    output n650;
    output n626;
    output n1381;
    output n904;
    output n1242;
    output n648;
    output n980;
    output n624;
    output n1382;
    output ootx_payloads_1_248;
    output ootx_payloads_1_247;
    output n902;
    output n1243;
    output n900;
    output n1244;
    output n978;
    output n674;
    output n1357;
    output n19;
    output n622;
    output n1383;
    output ootx_payloads_1_246;
    output ootx_payloads_1_245;
    output n898;
    output n1245;
    output ootx_payloads_1_244;
    output n896;
    output n1246;
    output n620;
    output n1384;
    output n6355;
    output n894;
    output n1247;
    output n6356;
    output n6357;
    output \ootx_payloads_N_1730[4] ;
    output n6358;
    output n750;
    output n1319;
    output n618;
    output n1385;
    output n892;
    output n1248;
    output n6359;
    output ootx_payloads_1_243;
    output n6361;
    output n890;
    output n1249;
    output ootx_payloads_1_242;
    output n6362;
    output n616;
    output n1386;
    output ootx_payloads_1_241;
    output ootx_payloads_1_240;
    output ootx_payloads_1_239;
    output n1006;
    output n888;
    output n1250;
    output ootx_payloads_1_238;
    output ootx_payloads_1_237;
    output n886;
    output n1251;
    output n614;
    output n1387;
    output n22943;
    output n976;
    output ootx_payloads_1_236;
    output n884;
    output n1252;
    output ootx_payloads_1_235;
    output n882;
    output n1253;
    output ootx_payloads_1_234;
    output n1358;
    output n612;
    output n1388;
    output n880;
    output n1254;
    output n748;
    output n1320;
    output n974;
    output n878;
    output n1255;
    output n1004;
    output n13329;
    output data_N_1808;
    output n6363;
    output n6364;
    output n6365;
    output ootx_payloads_1_233;
    input sensor_N_132;
    output n876;
    output n1256;
    output ootx_payloads_1_232;
    output n610;
    output n1389;
    output ootx_payloads_1_231;
    output n874;
    output n1257;
    output n872;
    output n1258;
    output n608;
    output n1390;
    output n870;
    output n1259;
    output n746;
    output n1321;
    output n606;
    output n1391;
    output n604;
    output n1392;
    output n710;
    output n1339;
    output n966;
    output n868;
    output n1260;
    output n602;
    output n1393;
    output n744;
    output n1322;
    output n866;
    output n1261;
    output n600;
    output n1394;
    output n864;
    output n1262;
    output n598;
    output n1395;
    output ootx_payloads_1_230;
    output ootx_payloads_1_229;
    output ootx_payloads_1_228;
    output ootx_payloads_1_227;
    output n596;
    output n1396;
    output n594;
    output n1397;
    output ootx_payloads_1_226;
    output ootx_payloads_1_225;
    output ootx_payloads_1_224;
    output n592;
    output n1398;
    output ootx_payloads_1_223;
    output n742;
    output n1323;
    output n862;
    output n1263;
    output n590;
    output n1399;
    output ootx_payloads_1_222;
    output ootx_payloads_1_221;
    output \ootx_payload_o[1][1] ;
    output ootx_payloads_1_220;
    output ootx_payloads_1_219;
    output ootx_payloads_1_218;
    output n588;
    output n1400;
    output ootx_payloads_1_217;
    output ootx_payloads_1_216;
    output \ootx_payload_o[1][2] ;
    output \ootx_payload_o[1][3] ;
    output \ootx_payload_o[1][4] ;
    output \ootx_payload_o[1][5] ;
    output \ootx_payload_o[1][6] ;
    output \ootx_payload_o[1][7] ;
    output \ootx_payload_o[1][8] ;
    output \ootx_payload_o[1][9] ;
    output \ootx_payload_o[1][10] ;
    output \ootx_payload_o[1][11] ;
    output \ootx_payload_o[1][12] ;
    output \ootx_payload_o[1][13] ;
    output \ootx_payload_o[1][14] ;
    output \ootx_payload_o[1][15] ;
    output \ootx_payload_o[1][16] ;
    output \ootx_payload_o[1][17] ;
    output \ootx_payload_o[1][18] ;
    output \ootx_payload_o[1][19] ;
    output \ootx_payload_o[1][20] ;
    output \ootx_payload_o[1][21] ;
    output \ootx_payload_o[1][22] ;
    output \ootx_payload_o[1][23] ;
    output \ootx_payload_o[1][24] ;
    output \ootx_payload_o[1][25] ;
    output \ootx_payload_o[1][26] ;
    output \ootx_payload_o[1][27] ;
    output \ootx_payload_o[1][28] ;
    output \ootx_payload_o[1][29] ;
    output \ootx_payload_o[1][30] ;
    output \ootx_payload_o[1][31] ;
    output \ootx_payload_o[1][32] ;
    output \ootx_payload_o[1][33] ;
    output \ootx_payload_o[1][34] ;
    output \ootx_payload_o[1][35] ;
    output \ootx_payload_o[1][36] ;
    output \ootx_payload_o[1][37] ;
    output \ootx_payload_o[1][38] ;
    output \ootx_payload_o[1][39] ;
    output \ootx_payload_o[1][40] ;
    output \ootx_payload_o[1][41] ;
    output \ootx_payload_o[1][42] ;
    output \ootx_payload_o[1][43] ;
    output \ootx_payload_o[1][44] ;
    output \ootx_payload_o[1][45] ;
    output \ootx_payload_o[1][46] ;
    output \ootx_payload_o[1][47] ;
    output \ootx_payload_o[1][48] ;
    output \ootx_payload_o[1][49] ;
    output \ootx_payload_o[1][50] ;
    output \ootx_payload_o[1][51] ;
    output \ootx_payload_o[1][52] ;
    output \ootx_payload_o[1][53] ;
    output \ootx_payload_o[1][54] ;
    output \ootx_payload_o[1][55] ;
    output \ootx_payload_o[1][56] ;
    output \ootx_payload_o[1][57] ;
    output \ootx_payload_o[1][58] ;
    output \ootx_payload_o[1][59] ;
    output \ootx_payload_o[1][60] ;
    output \ootx_payload_o[1][61] ;
    output \ootx_payload_o[1][62] ;
    output \ootx_payload_o[1][63] ;
    output \ootx_payload_o[1][64] ;
    output \ootx_payload_o[1][65] ;
    output \ootx_payload_o[1][66] ;
    output \ootx_payload_o[1][67] ;
    output \ootx_payload_o[1][68] ;
    output \ootx_payload_o[1][69] ;
    output \ootx_payload_o[1][70] ;
    output \ootx_payload_o[1][71] ;
    output \ootx_payload_o[1][72] ;
    output \ootx_payload_o[1][73] ;
    output \ootx_payload_o[1][74] ;
    output \ootx_payload_o[1][75] ;
    output \ootx_payload_o[1][76] ;
    output \ootx_payload_o[1][77] ;
    output \ootx_payload_o[1][78] ;
    output \ootx_payload_o[1][79] ;
    output \ootx_payload_o[1][80] ;
    output \ootx_payload_o[1][81] ;
    output \ootx_payload_o[1][82] ;
    output \ootx_payload_o[1][83] ;
    output \ootx_payload_o[1][84] ;
    output \ootx_payload_o[1][85] ;
    output \ootx_payload_o[1][86] ;
    output \ootx_payload_o[1][87] ;
    output \ootx_payload_o[1][88] ;
    output \ootx_payload_o[1][89] ;
    output \ootx_payload_o[1][90] ;
    output \ootx_payload_o[1][91] ;
    output \ootx_payload_o[1][92] ;
    output \ootx_payload_o[1][93] ;
    output \ootx_payload_o[1][94] ;
    output \ootx_payload_o[1][95] ;
    output \ootx_payload_o[1][96] ;
    output \ootx_payload_o[1][97] ;
    output \ootx_payload_o[1][98] ;
    output \ootx_payload_o[1][99] ;
    output \ootx_payload_o[1][100] ;
    output \ootx_payload_o[1][101] ;
    output \ootx_payload_o[1][102] ;
    output \ootx_payload_o[1][103] ;
    output \ootx_payload_o[1][104] ;
    output \ootx_payload_o[1][105] ;
    output \ootx_payload_o[1][106] ;
    output \ootx_payload_o[1][107] ;
    output \ootx_payload_o[1][108] ;
    output \ootx_payload_o[1][109] ;
    output \ootx_payload_o[1][110] ;
    output \ootx_payload_o[1][111] ;
    output \ootx_payload_o[1][112] ;
    output \ootx_payload_o[1][113] ;
    output \ootx_payload_o[1][114] ;
    output \ootx_payload_o[1][115] ;
    output \ootx_payload_o[1][116] ;
    output \ootx_payload_o[1][117] ;
    output \ootx_payload_o[1][118] ;
    output \ootx_payload_o[1][119] ;
    output \ootx_payload_o[1][120] ;
    output \ootx_payload_o[1][121] ;
    output \ootx_payload_o[1][122] ;
    output \ootx_payload_o[1][123] ;
    output \ootx_payload_o[1][124] ;
    output \ootx_payload_o[1][125] ;
    output \ootx_payload_o[1][126] ;
    output \ootx_payload_o[1][127] ;
    output \ootx_payload_o[1][128] ;
    output \ootx_payload_o[1][129] ;
    output \ootx_payload_o[1][130] ;
    output \ootx_payload_o[1][131] ;
    output \ootx_payload_o[1][132] ;
    output \ootx_payload_o[1][133] ;
    output \ootx_payload_o[1][134] ;
    output \ootx_payload_o[1][135] ;
    output \ootx_payload_o[1][136] ;
    output \ootx_payload_o[1][137] ;
    output \ootx_payload_o[1][138] ;
    output \ootx_payload_o[1][139] ;
    output \ootx_payload_o[1][140] ;
    output \ootx_payload_o[1][141] ;
    output \ootx_payload_o[1][142] ;
    output \ootx_payload_o[1][143] ;
    output \ootx_payload_o[1][144] ;
    output \ootx_payload_o[1][145] ;
    output \ootx_payload_o[1][146] ;
    output \ootx_payload_o[1][147] ;
    output \ootx_payload_o[1][148] ;
    output \ootx_payload_o[1][149] ;
    output \ootx_payload_o[1][150] ;
    output \ootx_payload_o[1][151] ;
    output \ootx_payload_o[1][152] ;
    output \ootx_payload_o[1][153] ;
    output \ootx_payload_o[1][154] ;
    output \ootx_payload_o[1][155] ;
    output \ootx_payload_o[1][156] ;
    output \ootx_payload_o[1][157] ;
    output \ootx_payload_o[1][158] ;
    output \ootx_payload_o[1][159] ;
    output \ootx_payload_o[1][160] ;
    output \ootx_payload_o[1][161] ;
    output \ootx_payload_o[1][162] ;
    output \ootx_payload_o[1][163] ;
    output \ootx_payload_o[1][164] ;
    output \ootx_payload_o[1][165] ;
    output \ootx_payload_o[1][166] ;
    output \ootx_payload_o[1][167] ;
    output \ootx_payload_o[1][168] ;
    output \ootx_payload_o[1][169] ;
    output \ootx_payload_o[1][170] ;
    output \ootx_payload_o[1][171] ;
    output \ootx_payload_o[1][172] ;
    output \ootx_payload_o[1][173] ;
    output \ootx_payload_o[1][174] ;
    output \ootx_payload_o[1][175] ;
    output \ootx_payload_o[1][176] ;
    output \ootx_payload_o[1][177] ;
    output \ootx_payload_o[1][178] ;
    output \ootx_payload_o[1][179] ;
    output \ootx_payload_o[1][180] ;
    output \ootx_payload_o[1][181] ;
    output \ootx_payload_o[1][182] ;
    output \ootx_payload_o[1][183] ;
    output \ootx_payload_o[1][184] ;
    output \ootx_payload_o[1][185] ;
    output \ootx_payload_o[1][186] ;
    output \ootx_payload_o[1][187] ;
    output \ootx_payload_o[1][188] ;
    output \ootx_payload_o[1][189] ;
    output \ootx_payload_o[1][190] ;
    output \ootx_payload_o[1][191] ;
    output \ootx_payload_o[1][192] ;
    output \ootx_payload_o[1][193] ;
    output \ootx_payload_o[1][194] ;
    output \ootx_payload_o[1][195] ;
    output \ootx_payload_o[1][196] ;
    output \ootx_payload_o[1][197] ;
    output \ootx_payload_o[1][198] ;
    output \ootx_payload_o[1][199] ;
    output \ootx_payload_o[1][200] ;
    output \ootx_payload_o[1][201] ;
    output \ootx_payload_o[1][202] ;
    output \ootx_payload_o[1][203] ;
    output \ootx_payload_o[1][204] ;
    output \ootx_payload_o[1][205] ;
    output \ootx_payload_o[1][206] ;
    output \ootx_payload_o[1][207] ;
    output \ootx_payload_o[1][208] ;
    output \ootx_payload_o[1][209] ;
    output \ootx_payload_o[1][210] ;
    output \ootx_payload_o[1][211] ;
    output \ootx_payload_o[1][212] ;
    output \ootx_payload_o[1][213] ;
    output \ootx_payload_o[1][214] ;
    output \ootx_payload_o[1][215] ;
    output \ootx_payload_o[1][216] ;
    output \ootx_payload_o[1][217] ;
    output \ootx_payload_o[1][218] ;
    output \ootx_payload_o[1][219] ;
    output \ootx_payload_o[1][220] ;
    output \ootx_payload_o[1][221] ;
    output \ootx_payload_o[1][222] ;
    output \ootx_payload_o[1][223] ;
    output \ootx_payload_o[1][224] ;
    output \ootx_payload_o[1][225] ;
    output \ootx_payload_o[1][226] ;
    output \ootx_payload_o[1][227] ;
    output \ootx_payload_o[1][228] ;
    output \ootx_payload_o[1][229] ;
    output \ootx_payload_o[1][230] ;
    output \ootx_payload_o[1][231] ;
    output \ootx_payload_o[1][232] ;
    output \ootx_payload_o[1][233] ;
    output \ootx_payload_o[1][234] ;
    output \ootx_payload_o[1][235] ;
    output \ootx_payload_o[1][236] ;
    output \ootx_payload_o[1][237] ;
    output \ootx_payload_o[1][238] ;
    output \ootx_payload_o[1][239] ;
    output \ootx_payload_o[1][240] ;
    output \ootx_payload_o[1][241] ;
    output \ootx_payload_o[1][242] ;
    output \ootx_payload_o[1][243] ;
    output \ootx_payload_o[1][244] ;
    output \ootx_payload_o[1][245] ;
    output \ootx_payload_o[1][246] ;
    output \ootx_payload_o[1][247] ;
    output \ootx_payload_o[1][248] ;
    output \ootx_payload_o[1][249] ;
    output \ootx_payload_o[1][250] ;
    output \ootx_payload_o[1][251] ;
    output \ootx_payload_o[1][252] ;
    output \ootx_payload_o[1][253] ;
    output \ootx_payload_o[1][254] ;
    output \ootx_payload_o[1][255] ;
    output \ootx_payload_o[1][256] ;
    output \ootx_payload_o[1][257] ;
    output \ootx_payload_o[1][258] ;
    output \ootx_payload_o[1][259] ;
    output \ootx_payload_o[1][260] ;
    output \ootx_payload_o[1][261] ;
    output \ootx_payload_o[1][262] ;
    output \ootx_payload_o[1][263] ;
    output n860;
    output n1264;
    output ootx_payloads_1_215;
    output n586;
    output n1401;
    output ootx_payloads_1_214;
    output n1359;
    output ootx_payloads_1_213;
    output ootx_payloads_1_212;
    output ootx_payloads_1_211;
    output n584;
    output n1402;
    output n582;
    output n1403;
    output ootx_payloads_1_210;
    output n858;
    output n1265;
    output ootx_payloads_1_209;
    output n580;
    output n1404;
    output ootx_payloads_1_208;
    output n578;
    output n1405;
    output n972;
    output n576;
    output n1406;
    output ootx_payloads_1_207;
    output ootx_payloads_1_206;
    output ootx_payloads_1_205;
    output ootx_payloads_1_204;
    output ootx_payloads_1_203;
    output n856;
    output n1266;
    output ootx_payloads_1_202;
    output n574;
    output n1407;
    output n970;
    output n968;
    output n572;
    output n1408;
    output ootx_payloads_1_201;
    output n854;
    output n1267;
    output n570;
    output n1409;
    output n740;
    output n1324;
    output ootx_payloads_1_200;
    output ootx_payloads_1_199;
    output n738;
    output n1325;
    output n568;
    output n1410;
    output ootx_payloads_1_198;
    output n852;
    output n1268;
    output ootx_payloads_1_197;
    output n566;
    output n1411;
    output ootx_payloads_1_196;
    output ootx_payloads_1_195;
    output ootx_payloads_1_194;
    output ootx_payloads_1_193;
    output ootx_payloads_1_192;
    output n564;
    output n1412;
    output n850;
    output n1269;
    output n1360;
    output n562;
    output n1413;
    output n708;
    output n1340;
    output n560;
    output n1414;
    output n964;
    output n9513;
    input ootx_payloads_N_1698;
    output n558;
    output n1415;
    output ootx_payloads_1_191;
    output ootx_payloads_1_190;
    output ootx_payloads_1_189;
    output ootx_payloads_1_188;
    output ootx_payloads_1_187;
    output n848;
    output n1270;
    output ootx_payloads_1_186;
    output n556;
    output n1416;
    output ootx_payloads_1_185;
    output ootx_payloads_1_184;
    output n554;
    output n1417;
    output ootx_payloads_1_183;
    output n768;
    output n1310;
    output n846;
    output n1271;
    output ootx_payloads_1_182;
    output n540;
    output n542;
    output n544;
    output n546;
    output n548;
    output ootx_payloads_1_181;
    output n550;
    output n552;
    output n1370;
    output n736;
    output n686;
    output n690;
    output ootx_payloads_1_180;
    output n762;
    output n692;
    output ootx_payloads_1_179;
    output n1313;
    output n696;
    output n698;
    output ootx_payloads_1_178;
    output n700;
    output n702;
    output ootx_payloads_1_177;
    output n936;
    output n1226;
    output ootx_payloads_1_176;
    output n704;
    output ootx_payloads_1_175;
    output ootx_payloads_1_174;
    output n706;
    output ootx_payloads_1_173;
    output ootx_payloads_1_172;
    output ootx_payloads_1_171;
    output ootx_payloads_1_170;
    output ootx_payloads_1_169;
    output ootx_payloads_1_168;
    output ootx_payloads_1_167;
    output ootx_payloads_1_166;
    output ootx_payloads_1_165;
    output n962;
    output ootx_payloads_1_164;
    output ootx_payloads_1_163;
    output ootx_payloads_1_162;
    output n646;
    output n1371;
    output ootx_payloads_1_161;
    output ootx_payloads_1_160;
    output n720;
    output ootx_payloads_1_159;
    output n760;
    output ootx_payloads_1_158;
    output n1314;
    output n642;
    output n644;
    output ootx_payloads_1_157;
    output ootx_payloads_1_156;
    output ootx_payloads_1_155;
    output ootx_payloads_1_154;
    output ootx_payloads_1_153;
    output ootx_payloads_1_152;
    output ootx_payloads_1_151;
    output ootx_payloads_1_150;
    output ootx_payloads_1_149;
    output ootx_payloads_1_148;
    output ootx_payloads_1_147;
    output n960;
    output ootx_payloads_1_146;
    output n770;
    output n772;
    output ootx_payloads_1_145;
    output n774;
    output n718;
    output ootx_payloads_1_144;
    output ootx_payloads_1_143;
    output n1361;
    output n682;
    output n684;
    output ootx_payloads_1_142;
    output n688;
    output ootx_payloads_1_141;
    output ootx_payloads_1_140;
    output n694;
    output ootx_payloads_1_139;
    output ootx_payloads_1_138;
    output ootx_payloads_1_137;
    output ootx_payloads_1_136;
    output ootx_payloads_1_135;
    output n734;
    output n776;
    output ootx_payloads_1_134;
    output ootx_payloads_1_133;
    output ootx_payloads_1_132;
    output ootx_payloads_1_131;
    output n538;
    output n756;
    output n758;
    output ootx_payloads_1_130;
    output ootx_payloads_1_129;
    output n728;
    output ootx_payloads_1_128;
    output ootx_payloads_1_127;
    output n714;
    output n730;
    output n732;
    output ootx_payloads_1_126;
    output ootx_payloads_1_125;
    output ootx_payloads_1_124;
    output ootx_payloads_1_123;
    output ootx_payloads_1_122;
    output n716;
    output ootx_payloads_1_121;
    output ootx_payloads_1_120;
    output ootx_payloads_1_119;
    output ootx_payloads_1_118;
    output ootx_payloads_1_117;
    output ootx_payloads_1_116;
    output ootx_payloads_1_115;
    output n1315;
    output ootx_payloads_1_114;
    output n722;
    output ootx_payloads_1_113;
    output ootx_payloads_1_112;
    output ootx_payloads_1_111;
    output n1333;
    output ootx_payloads_1_110;
    output n726;
    output ootx_payloads_1_109;
    output ootx_payloads_1_108;
    output ootx_payloads_1_107;
    output n1418;
    output ootx_payloads_1_106;
    output ootx_payloads_1_105;
    output ootx_payloads_1_104;
    output ootx_payloads_1_103;
    output ootx_payloads_1_102;
    output ootx_payloads_1_101;
    output n1216;
    output n844;
    output n1272;
    output n1217;
    output ootx_payloads_1_100;
    output n1218;
    output ootx_payloads_1_99;
    output n1219;
    output n842;
    output n1273;
    output n1419;
    output n1220;
    output ootx_payloads_1_98;
    output ootx_payloads_1_97;
    output ootx_payloads_1_96;
    output n1221;
    output ootx_payloads_1_95;
    output ootx_payloads_1_94;
    output ootx_payloads_1_93;
    output n1222;
    output ootx_payloads_1_92;
    output n1341;
    output ootx_payloads_1_91;
    output n1223;
    output ootx_payloads_1_90;
    output n1224;
    output ootx_payloads_1_89;
    output ootx_payloads_1_88;
    output ootx_payloads_1_87;
    output ootx_payloads_1_86;
    output n840;
    output n1274;
    output ootx_payloads_1_85;
    output ootx_payloads_1_84;
    output ootx_payloads_1_83;
    output n1420;
    output n1227;
    output ootx_payloads_1_82;
    output n1228;
    output n838;
    output n1275;
    output ootx_payloads_1_81;
    output n934;
    output n1229;
    output ootx_payloads_1_80;
    output ootx_payloads_1_79;
    output ootx_payloads_1_78;
    output ootx_payloads_1_77;
    output ootx_payloads_1_76;
    output ootx_payloads_1_75;
    output n1342;
    output n1421;
    output ootx_payloads_1_74;
    output n836;
    output n1276;
    output ootx_payloads_1_73;
    output ootx_payloads_1_72;
    output n1422;
    output n1423;
    output n834;
    output n1277;
    output ootx_payloads_1_71;
    output ootx_payloads_1_70;
    output n1424;
    output ootx_payloads_1_69;
    output ootx_payloads_1_68;
    output ootx_payloads_1_67;
    output ootx_payloads_1_66;
    output ootx_payloads_1_65;
    output ootx_payloads_1_64;
    output n1343;
    output n1425;
    output ootx_payloads_1_63;
    output n832;
    output n1278;
    output ootx_payloads_1_62;
    output ootx_payloads_1_61;
    output n536;
    output n1426;
    output n1316;
    output ootx_payloads_1_60;
    output n1334;
    output ootx_payloads_1_59;
    output ootx_payloads_1_58;
    output ootx_payloads_1_57;
    output n534;
    output n1427;
    output ootx_payloads_1_56;
    output n830;
    output n1279;
    output n1362;
    output ootx_payloads_1_55;
    output ootx_payloads_1_54;
    output ootx_payloads_1_53;
    output n1344;
    output n532;
    output n1428;
    output ootx_payloads_1_52;
    output n828;
    output n1280;
    output n530;
    output n1429;
    output n956;
    output n1345;
    output ootx_payloads_1_51;
    output ootx_payloads_1_50;
    output ootx_payloads_1_49;
    output n954;
    output n826;
    output n1281;
    output ootx_payloads_1_48;
    output n528;
    output n1430;
    output ootx_payloads_1_47;
    output n526;
    output n1431;
    output ootx_payloads_1_46;
    output ootx_payloads_1_45;
    output n1346;
    output n824;
    output n1282;
    output ootx_payloads_1_44;
    output n952;
    output ootx_payloads_1_43;
    output n524;
    output n1432;
    output \ootx_payloads_N_1730[12] ;
    output ootx_payloads_1_42;
    output ootx_payloads_1_41;
    output ootx_payloads_1_40;
    output ootx_payloads_1_39;
    output ootx_payloads_1_38;
    output ootx_payloads_1_37;
    output n522;
    output n1433;
    output n822;
    output n1283;
    output n1347;
    output n950;
    output \ootx_payloads_N_1730[11] ;
    output ootx_payloads_1_36;
    output ootx_payloads_1_35;
    output n1326;
    output ootx_payloads_1_34;
    output ootx_payloads_1_33;
    output n1348;
    output n6334;
    output ootx_payloads_1_32;
    output ootx_payloads_1_31;
    output n51;
    output n52;
    output ootx_payloads_1_30;
    output n948;
    output \ootx_payloads_N_1730[10] ;
    output ootx_payloads_1_29;
    output ootx_payloads_1_28;
    input n2679;
    input n2680;
    output n6335;
    output n1349;
    output ootx_payloads_1_27;
    output n1317;
    output n932;
    output ootx_payloads_1_26;
    output n6336;
    output n946;
    output ootx_payloads_1_25;
    output ootx_payloads_1_24;
    output ootx_payloads_1_23;
    output \ootx_payloads_N_1730[9] ;
    output n1363;
    output ootx_payloads_1_22;
    output n49;
    output n50;
    output n9771;
    output n820;
    output n1284;
    output ootx_payloads_1_21;
    output n6337;
    output ootx_payloads_1_20;
    output n1350;
    output ootx_payloads_1_19;
    output ootx_payloads_1_18;
    output ootx_payloads_1_17;
    output n944;
    output n6338;
    output ootx_payloads_1_16;
    output n1351;
    output \ootx_payloads_N_1730[8] ;
    output n47;
    output n48;
    output n818;
    output n1285;
    output ootx_payloads_1_15;
    output ootx_payloads_1_14;
    output ootx_payloads_1_13;
    output ootx_payloads_1_12;
    output n942;
    output n6339;
    output ootx_payloads_1_11;
    output n45;
    output n46;
    output ootx_payloads_1_10;
    output \ootx_payloads_N_1730[7] ;
    output n816;
    output n1286;
    output ootx_payloads_1_9;
    output n6340;
    output ootx_payloads_1_8;
    output crc32s_1_25;
    output crc32s_1_30;
    output crc32s_1_27;
    output crc32s_1_26;
    output crc32s_1_31;
    output crc32s_1_29;
    output crc32s_1_28;
    output crc32s_1_24;
    output crc32s_1_23;
    output crc32s_1_22;
    output crc32s_1_21;
    output ootx_payloads_1_7;
    output crc32s_1_20;
    output \ootx_payloads_N_1730[6] ;
    output n1364;
    output ootx_payloads_1_6;
    output ootx_payloads_1_5;
    output crc32s_1_19;
    output crc32s_1_18;
    output crc32s_1_17;
    output crc32s_1_16;
    output crc32s_1_15;
    output n6341;
    output crc32s_1_14;
    output crc32s_1_13;
    output crc32s_1_12;
    output crc32s_1_11;
    output crc32s_1_10;
    output crc32s_1_9;
    output crc32s_1_8;
    output crc32s_1_7;
    output crc32s_1_6;
    output crc32s_1_5;
    output crc32s_1_4;
    output crc32s_1_3;
    output crc32s_1_2;
    output ootx_payloads_1_4;
    output ootx_payloads_1_3;
    output crc32s_1_0;
    output ootx_payloads_1_2;
    output crc32s_1_1;
    output \ootx_payloads_N_1730[5] ;
    output ootx_payloads_1_1;
    output n43;
    output n6342;
    output n44;
    output n28;
    output n814;
    output n1287;
    output n41;
    output n42;
    output n1288;
    output n1289;
    output n1290;
    output n1291;
    output n1292;
    output n1293;
    output n1294;
    output n1295;
    output n1296;
    output n1297;
    output n1298;
    output n1299;
    output n1300;
    output n1301;
    output n1302;
    output n1303;
    output n1304;
    output n1305;
    output n1306;
    output n1307;
    output n1308;
    output n1309;
    output n1327;
    output n1328;
    output n1329;
    output n1330;
    output n1331;
    output n1335;
    output n1336;
    output n1337;
    output n1352;
    output n1353;
    output n1365;
    output n1366;
    output n1367;
    output n1368;
    output n1369;
    output n1372;
    output n1373;
    input n11612;
    output [31:0]n3112;
    input n11611;
    input n11610;
    input n11609;
    input n11608;
    input n11607;
    input n11606;
    input n11605;
    input n11604;
    input n22997;
    input n11602;
    input n23001;
    input n11600;
    input n11599;
    input n11598;
    input n11597;
    input n11596;
    input n11595;
    input n11594;
    input n11593;
    input n11592;
    input n11591;
    input n11590;
    input n11589;
    input n11588;
    input n11587;
    input n11586;
    input n11585;
    input n11584;
    input n11583;
    input n11582;
    input n11581;
    input n11580;
    input n11579;
    input n11578;
    input n11577;
    input n11576;
    input n11575;
    input n11574;
    input n11573;
    input n11572;
    input n11571;
    input n11570;
    input n11569;
    input n11568;
    input n11567;
    input n11566;
    input n11565;
    input n11564;
    input n11563;
    input n11562;
    input n11561;
    input n11560;
    input n11559;
    input n11558;
    input n11557;
    input n11556;
    input n11555;
    input n11554;
    input n11553;
    input n11552;
    input n11551;
    input n11550;
    input n11549;
    input n11548;
    input n11547;
    input n11546;
    input n11545;
    input n11544;
    input n11543;
    input n11542;
    input n11541;
    input n11540;
    input n11539;
    input n11538;
    input n11537;
    input n11536;
    input n11535;
    input n11534;
    input n11533;
    input n11532;
    input n11531;
    input n11530;
    input n11529;
    input n11528;
    input n11527;
    input n11526;
    input n11525;
    input n11524;
    input n11523;
    input n11522;
    input n11521;
    input n11520;
    input n11519;
    input n11518;
    input n11517;
    input n11516;
    input n11515;
    input n11514;
    input n11513;
    input n11512;
    input n11511;
    input n11510;
    input n11509;
    input n11508;
    input n11507;
    input n11506;
    input n11505;
    input n11504;
    output n39;
    output n40;
    output n812;
    output n37;
    output n38;
    output n6343;
    output n810;
    output n808;
    output n17;
    output n19468;
    output n806;
    output n535;
    output n792;
    output n804;
    output n533;
    output led_c_0;
    output n790;
    output led_c_1;
    output led_c_2;
    output led_c_3;
    output led_c_4;
    output led_c_5;
    output led_c_6;
    output n802;
    output n800;
    output n531;
    input n11503;
    input n11502;
    input n11501;
    input n11500;
    input n11499;
    input n11498;
    input n11497;
    input n11496;
    input n11495;
    input n11494;
    input n11493;
    input n11492;
    input n11491;
    input n11490;
    input n11489;
    input n11488;
    input n11487;
    input n11486;
    input n11485;
    input n11484;
    input n11483;
    input n11482;
    input n11481;
    input n11480;
    input n11479;
    input n11478;
    input n11477;
    input n11476;
    input n11475;
    input n11474;
    input n11473;
    input n11472;
    output n788;
    input n11471;
    input n11470;
    input n11469;
    input n11468;
    input n11467;
    input n11466;
    input n11465;
    input n11464;
    input n11463;
    input n11462;
    input n11461;
    input n11460;
    input n11459;
    input n11458;
    input n11457;
    input n11456;
    input n11455;
    input n11454;
    input n11453;
    input n11452;
    input n11451;
    input n11450;
    input n11449;
    input n11448;
    input n11447;
    input n11446;
    input n11445;
    input n11444;
    input n11443;
    input n11442;
    input n11441;
    input n11440;
    input n11439;
    input n11438;
    input n11437;
    input n11436;
    input n11435;
    input n11434;
    input n11433;
    input n11432;
    input n11431;
    input n11430;
    input n11429;
    input n11428;
    input n11427;
    input n11426;
    input n11425;
    input n11424;
    input n11423;
    input n11422;
    input n11421;
    input n11420;
    input n11419;
    input n11418;
    input n11417;
    input n11416;
    input n11415;
    input n11414;
    input n11413;
    input n11412;
    input n11411;
    input n11410;
    input n11409;
    input n11408;
    input n11407;
    input n11406;
    input n11405;
    input n11404;
    input n11403;
    input n11402;
    input n11401;
    input n11400;
    input n11399;
    input n11398;
    input n11397;
    input n11396;
    input n11395;
    input n11394;
    input n11393;
    input n11392;
    input n11391;
    input n11390;
    input n11389;
    input n11388;
    input n11387;
    input n11386;
    input n11385;
    input n11384;
    input n11383;
    input n11382;
    input n11381;
    input n11380;
    input n11379;
    input n11378;
    input n11377;
    input n11376;
    input n11375;
    input n11374;
    input n11373;
    input n11372;
    input n11371;
    input n11370;
    input n11369;
    input n11368;
    input n11367;
    input n11366;
    input n11365;
    input n11364;
    input n11363;
    input n11362;
    input n11361;
    input n11360;
    input n11359;
    input n11358;
    input n11357;
    input n11356;
    input n11355;
    input n11354;
    input n11353;
    input n11352;
    input n11351;
    input n11350;
    input n11349;
    input n11348;
    input n11347;
    input n11346;
    input n11345;
    input n11344;
    input n11343;
    input n11342;
    input n11341;
    input n11340;
    input n11339;
    input n11338;
    input n11337;
    input n11336;
    input n11335;
    input n11334;
    input n11333;
    input n11332;
    input n11331;
    input n11330;
    input n11329;
    input n11328;
    input n11327;
    input n11326;
    input n11325;
    input n11324;
    input n11323;
    input n11322;
    input n11321;
    input n11320;
    input n11319;
    input n11318;
    input n11317;
    input n11316;
    input n11315;
    input n11314;
    input n11313;
    input n11312;
    input n11311;
    input n11310;
    input n11309;
    input n11308;
    input n11307;
    input n11306;
    input n11305;
    input n11304;
    input n11303;
    input n11302;
    input n11301;
    input n11300;
    input n11299;
    input n11298;
    input n11297;
    input n11296;
    input n11295;
    input n11294;
    input n11293;
    input n11292;
    input n11291;
    input n11290;
    input n11289;
    input n11288;
    input n11287;
    input n11286;
    input n11285;
    output ootx_payloads_1_0;
    output n6344;
    output n798;
    output n529;
    output n796;
    output n6345;
    output n786;
    output n794;
    output n527;
    output n6346;
    output n784;
    output n525;
    output n782;
    output n523;
    output n780;
    output n778;
    output n521;
    output n1032;
    output \ootx_payloads_N_1730[0] ;
    output n930;
    output n940;
    output [1:0]sync;
    output n1022;
    output n1012;
    output n1014;
    output n1002;
    output n1016;
    output n1018;
    output n1020;
    output n1024;
    output n1026;
    output n1028;
    output n1030;
    input n11016;
    output \ootx_payload_o[0][0] ;
    output n67;
    output n65;
    output n63;
    output \ootx_states[1][0] ;
    input n25;
    output n61;
    output n59;
    output n57;
    output n55;
    output n53;
    output n68;
    output n66;
    output n64;
    output n62;
    output n60;
    output n58;
    output n56;
    output n54;
    input n20_adj_33;
    output led_c_7;
    
    wire clock_c /* synthesis SET_AS_NETWORK=clock_c, is_clock=1 */ ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/DarkRoomOOTXdecoder.v(40[8:13])
    
    wire ootx_shift_registers_N_1748, ootx_shift_registers_1_3, ootx_shift_registers_1_4, 
        n11045, n2297, n2198, n2225, n22601, n22292, n3017, n25183;
    wire [271:0]n2;
    
    wire n2283, n22477, n1503, n1532, n22478, n2891, n2792, n2819, 
        n22748, n2691, n2592, n2621, n22697, n22698, n22602, n22293, 
        n2324, n25198, ootx_shift_registers_1_1, ootx_shift_registers_1_2, 
        n11043, n22291, n1119, crc32s_N_1751, n10243, n22972, n1087, 
        n1603, n1504, n22476, n22749, n11852, payload_lengths_0_1, 
        payload_lengths_1_1, n2298, n2199, n22600, n2692, n2593, 
        n22696, n3212, n25181, n22812, ootx_shift_registers_1_0, n11041, 
        n1604, n1505, n22475, n2299, n2200, n22599;
    wire [30:0]n2849;
    
    wire n22261, n2984, n2885, n2918, n22782, ootx_payloads_0_239, 
        n11260, n22262, n2892, n2793, n22747, n2693, n2594, n22695, 
        n22813, n11044, n1605, n1506, n22474, n11144, ootx_payloads_0_123, 
        n2093, n2099, n2103, n26, n2098, n2104, n2097, n2105, 
        n29, n2300, n2201, n22598, n22290, n2112, n2111, n2110, 
        n22941, n11143, ootx_payloads_0_122, n2096, n2102, n20_c, 
        payload_lengths_0_2, payload_lengths_1_2, n2100, n2101, n2108, 
        n2107, n28_c, n2095, n2106, n32, n11142, ootx_payloads_0_121, 
        n2985, n2886, n22781;
    wire [30:0]ootx_payloads_N_1699;
    
    wire n8941, n88, n17_c, n11141, ootx_payloads_0_120, n20112, 
        n11140, ootx_payloads_0_119, n1712, n1711, n1710, n22946, 
        n11139, ootx_payloads_0_118, n1699, n1706_adj_1810, n16, n2094, 
        n2109, n19_c, n1704, n1707, n1700, n1701, n22, n11138, 
        ootx_payloads_0_117, n2126, n1705, n1709, n1702, n20_adj_1811, 
        n1697, n1708, n24, n11137, ootx_payloads_0_116, n20105, 
        n11136, ootx_payloads_0_115, n23985, n1698, n1703, n1730, 
        n11135, ootx_payloads_0_114, n11134, ootx_payloads_0_113, n1606, 
        n1507, n22473, n22260, n2720, n25192, n11133, ootx_payloads_0_112, 
        n11132, ootx_payloads_0_111, payload_lengths_0_3, payload_lengths_1_3, 
        n11131, ootx_payloads_0_110, n11130, ootx_payloads_0_109, n2301, 
        n2202, n22597, n22231, n4, n11129, ootx_payloads_0_108, 
        n11128, ootx_payloads_0_107;
    wire [30:0]n69;
    
    wire n11127, ootx_payloads_0_106, n2986, n2887, n22780, n11126, 
        ootx_payloads_0_105, n22232, n11851, ootx_payloads_0_238, n11259, 
        n11125, ootx_payloads_0_104, n11850, n2694, n2595, n22694, 
        n25182, ootx_payloads_0_237, n11258, n1607, n1508, n22472, 
        n22259, n11849, n2302, n2203, n22596, n2695, n2596, n22693, 
        n1608, n1509, n25177, n22471, n22289, ootx_payloads_0_236, 
        n11257, n2303, n2204, n22595, n22258, n11848, n22230, 
        n2987, n2888, n22779, n3083, n22811, ootx_payloads_0_235, 
        n11256, n2893, n2794, n22746, n2988, n2889, n22778, n11735, 
        n9498, n118, n11847, n1609, n1510, n22470, ootx_payloads_0_234, 
        n11255, n2304, n2205, n22594, n2696, n2597, n22692, n1829, 
        n25196;
    wire [31:0]n71;
    
    wire n839, n912_c, n1812, n1811, n1810, n22945, n1610, n1511, 
        n22469, n22288, n2305, n2206, n22593, n2697, n2598, n22691, 
        n11846, n1799, n1809, n18, ootx_payloads_0_233, n11254, 
        n1805, n1802, n1803, n1797, n24_adj_1812, n1807, n1796, 
        n1806, n1800, n22_adj_1813, n2894, n2795, n22745;
    wire [1:0]n72;
    
    wire n1808, n1801, n26_adj_1815, n1804, n1798, n22287, n1611, 
        n1512, n22468, n24028, n24829, n11124, ootx_payloads_0_103, 
        n3084, n22810, n2306, n2207, n22592, n11123, ootx_payloads_0_102, 
        n811, n910_c, n938_c, n25195, n11122, ootx_payloads_0_101, 
        n11121, ootx_payloads_0_100, n11120, ootx_payloads_0_99, n2698, 
        n2599, n22690, n10357, n809, n908_c, n808_c, n907, n2895, 
        n2796, n22744, n1928, n25191, n22257, n807, n906_c;
    wire [31:0]n773;
    
    wire n740_c, n812_c, n711, n810_c, n1612, n909, n911, n11845, 
        n709, n708_c, ootx_payloads_0_232, n11253, n27, n712_c, 
        n58_c, n24097, n3085, n22809, n610_c;
    wire [31:0]n89;
    
    wire n641, n62_c, n24124, n2307, n2208, n22591, n66_c, n24095, 
        n70, n24093, payload_lengths_0_4, n74, n24091, payload_lengths_0_5, 
        n11119, ootx_payloads_0_98, n78, n24089, payload_lengths_0_6, 
        n82, n24087, payload_lengths_0_7, n86, n24085, payload_lengths_0_8, 
        n90, n24083, payload_lengths_0_9, n94, n24081, payload_lengths_0_10, 
        n98, n24079, payload_lengths_0_11, n102, n24077, payload_lengths_0_12, 
        n106, n24075, payload_lengths_0_13, n11118, ootx_payloads_0_97, 
        n110, n24073, payload_lengths_0_14, n114, n24071, payload_lengths_0_15, 
        n122, n24069, n609, n126, n24067, n58_adj_1820, n60_c, 
        n130, n24065, n134, n24063, payload_lengths_1_4, n138, n24061, 
        payload_lengths_1_5, n11117, ootx_payloads_0_96, n142, n24059, 
        payload_lengths_1_6, n146, n24057, payload_lengths_1_7, n150, 
        n24055, payload_lengths_1_8, n154, n24053, payload_lengths_1_9, 
        n158, n24051, payload_lengths_1_10, n162, n24049, payload_lengths_1_11, 
        n166, n24047, payload_lengths_1_12, n170, n24045, payload_lengths_1_13, 
        n11116, ootx_payloads_0_95;
    wire [31:0]n91;
    wire [31:0]counter_from_nskip_rise;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(36[9:32])
    
    wire n174, n24043, payload_lengths_1_14, n178, n24041, payload_lengths_1_15, 
        n23689;
    wire [31:0]counter_from_last_rise_c;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    
    wire n11844;
    wire [1:0]ootx_states_1__1__N_896;
    
    wire n23147;
    wire [1:0]\ootx_states[1] ;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(52[9:20])
    
    wire n11115, ootx_payloads_0_94, n31, n22_adj_1846, n34_c, ootx_payloads_0_231, 
        n11252, n11821, n83, n19313, n608_c, n23163, n2989, n2890, 
        n22777, n22286, n22256, n11831, n2699, n2600, n22689, 
        n22229, n10802;
    wire [1:0]ootx_states_0__1__N_898;
    
    wire ootx_payloads_0_218, n11239, n1499, n1400_c, n1433_c, n22467, 
        n2308, n2209, n25179, n22590, n1500, n1401_c, n22466, 
        n2700, n2601, n22688, n11843, ootx_payloads_0_230, n11251, 
        n11114, ootx_payloads_0_93, ootx_payloads_0_208, n11229, n612_c, 
        n611, n22887, n2309, n2210, n22589, n1501, n1402_c, n22465, 
        n2896, n2797, n22743, n22255, n2701, n2602, n22687, n23693, 
        n22285, n710_c, n22886, n707, n22254, n11113, ootx_payloads_0_92, 
        ootx_payloads_0_79, n11100, n11692, n806_c, n23950, n6, 
        n29_adj_1850, n11708, n24713, n24553, n4_adj_1851, n39_c, 
        n905, n29_adj_1852, n126_adj_1853, n125, n13_adj_1854, n30_adj_1855, 
        n1037, n25193, n2412, n2411, n2410, n22896, n2408, n2409, 
        n23, n2404, n2403, n2407, n2398, n31_adj_1856, n24697;
    wire [31:0]n6333_c;
    
    wire n2399, n2392, n36, n2391, n2394, n2393, n2402, n34_adj_1857, 
        n2390, n2400, n2396, n2405, n35_adj_1858, n2406, n2397, 
        n2395, n2401, n33, n22228, n3086, n22808, n2423, n1005, 
        n1006_c, n1008_c, n1004_c, n10;
    wire [14:0]n4485;
    
    wire n1012_c, n1011, n1010_c, n22876, n1007, n1009, n11112, 
        ootx_payloads_0_91, n11111, ootx_payloads_0_90, n11110, ootx_payloads_0_89, 
        n11109, ootx_payloads_0_88, n11108, ootx_payloads_0_87, n11107, 
        ootx_payloads_0_86, n38_c, n86_adj_1860, n85, n11106, ootx_payloads_0_85, 
        n2310, n2211, n22588, n11105, ootx_payloads_0_84, n11104, 
        ootx_payloads_0_83, ootx_payloads_N_1685, n11103, ootx_payloads_0_82, 
        n1502, n1403_c, n22464, n1912, n1911, n1910, n22944, n1906, 
        n1900, n1903, n1905, n26_adj_1861, n11938, n11937, n11936, 
        n11935, n11934, n11933, n11932, n11931, n11930, n11929, 
        n11928, n11927, n11926, n1898, n1895, n1896, n1897, n24_adj_1862, 
        n1904, n1902, n1901, n1899, n25_c, n1908, n1909, n1907, 
        n23_adj_1863, n2522, n25187, n1136, n25190, n11925, n11924, 
        n11923, n11922, n11921, n11920, n11919, n11918, n11917, 
        n11916, n11915, n11914, n11913, n11912, n11911, n11910, 
        n11909, n11908, n11907, n11906, n11905, n11904, n11903, 
        n11902, n11901, n11900, n11899, n17_adj_1864, n18_adj_1865, 
        n11898, n11897, n11896, n11895, n11894, n11893, n11892, 
        n11891, n11890, n11889, n11888, n11887, n11886, n11885, 
        n11884, n11883, n11882, n11881, n11880, n11879, n11878, 
        n11877, n11876, n11875, n11874, n11873, n11872, n11871, 
        n11870, n11869, n11868, n2712, n2711, n2710, n22893, n11867, 
        n2690, n2708, n2689, n36_adj_1866, n11866, n11865, n11864, 
        n11863, n11862, n2703, n2709, n32_adj_1867, n11861, n11860, 
        n2706, n2707, n2704, n2705, n40_c, n11859, n11858, n2688, 
        n38_adj_1868, n11857, n11856, n11102, ootx_payloads_0_81, 
        n2702, n37_c, n2687, n41_c, n43_adj_1869, n2027, n25188, 
        n2311, n2212, n22587, n11855, n11854, n1404_c, n22463, 
        n2990, n22776, n11853, n11101, ootx_payloads_0_80, n1108, 
        n1103, n8_adj_1870, n1106, n1107, n1104, n1105, n12, n1112, 
        n1111, n1110, n22906, n11672, n3087, n22807, ootx_payloads_0_59, 
        n11080, n11816, n2991, n22775, n11842, n11841, n2897, 
        n2798, n22742, n11840, n11839, n11838, n1109, n11837, 
        n11836, n11714, n2603, n22686, n1235_c, n25189, n11835, 
        n11834, ootx_payloads_0_203, n11224, n11833, n113, n11832, 
        n96, n11671, ootx_payloads_0_263, ootx_payloads_0_58, n11079, 
        n11815, ootx_payloads_0_202, n11223, n94_adj_1872, n82_adj_1873, 
        n432, n11734, n23_adj_1874, ootx_payloads_0_262, n81, n11814, 
        ootx_payloads_0_201, n11222, n11670, ootx_payloads_0_57, n11078, 
        n92, n11813, ootx_payloads_0_200, n11221, n11669, ootx_payloads_0_56, 
        n11077, n90_adj_1876, n11812, ootx_payloads_0_199, n11220, 
        n11668, ootx_payloads_0_55, n11076, n88_adj_1877, n11811, 
        ootx_payloads_0_198, n11219, n11810, ootx_payloads_0_197, n11218, 
        n11728, n84, n11809, ootx_payloads_0_196, n11217, n4729, 
        n11691, n11808, ootx_payloads_0_195, n11216, ootx_shift_registers_0_13, 
        ootx_shift_registers_1_13;
    wire [17:0]data_counters_N_1780;
    
    wire ootx_shift_registers_0_0, ootx_shift_registers_0_14, ootx_shift_registers_1_14, 
        ootx_shift_registers_0_6, ootx_shift_registers_1_6, ootx_shift_registers_0_9, 
        ootx_shift_registers_1_9, ootx_shift_registers_0_15, ootx_shift_registers_1_15, 
        ootx_shift_registers_0_10, ootx_shift_registers_1_10, n20_adj_1881, 
        ootx_shift_registers_0_4, ootx_shift_registers_0_2, n19_adj_1882, 
        ootx_shift_registers_0_17, ootx_shift_registers_1_17, ootx_shift_registers_0_7, 
        ootx_shift_registers_1_7, ootx_shift_registers_0_16, ootx_shift_registers_1_16, 
        ootx_shift_registers_0_11, ootx_shift_registers_1_11, n24_adj_1883, 
        ootx_shift_registers_0_12, ootx_shift_registers_1_12, n22_adj_1884, 
        ootx_shift_registers_0_5, ootx_shift_registers_1_5, n23_adj_1885, 
        n11667, ootx_payloads_0_261, ootx_payloads_0_54, n11075, ootx_payloads_0_260, 
        ootx_payloads_0_78, n11099, n80, ootx_payloads_0_259, n3088, 
        n22806, n11807, ootx_shift_registers_0_1, n21, ootx_shift_registers_0_3, 
        n26_adj_1887, n32_adj_1888, ootx_shift_registers_0_8, ootx_shift_registers_1_8, 
        n25_adj_1889, n33_adj_1890, ootx_payloads_0_194, n11215, n24133, 
        data_counters_N_1776, n78_adj_1891, n111, n11690, n11806, 
        ootx_payloads_0_258, n2992, n22774, ootx_payloads_0_193, n11214, 
        ootx_payloads_0_257, ootx_payloads_0_256, n11666, ootx_payloads_0_255, 
        n10_adj_1895, n16_adj_1896, n15, n4_adj_1897, ootx_payloads_0_254, 
        ootx_payloads_0_53, n11074, ootx_payloads_0_253, n76, ootx_payloads_0_252, 
        n23741, ootx_payloads_0_77, n11098, ootx_payloads_0_251, n11805, 
        ootx_payloads_0_250, ootx_payloads_0_249, ootx_payloads_0_192, 
        n11213, n74_adj_1899, n14, n13_adj_1900, n15_adj_1901, n24013, 
        n11665, ootx_payloads_0_52, n11073, n11804, ootx_payloads_0_191, 
        n11212, n39_adj_1902, n135, n24_adj_1903, n79, n136, n11664, 
        ootx_payloads_0_248, ootx_payloads_0_229, n11250, ootx_payloads_0_51, 
        n11072, ootx_payloads_0_247, n11803, ootx_payloads_0_190, n11211, 
        n11802, ootx_payloads_0_189, n11210, n66_adj_1904, n162_adj_1905, 
        ootx_payloads_0_228, n11249, n11689, n11663, ootx_payloads_0_246, 
        ootx_payloads_0_245, ootx_payloads_0_50, n11071, n11801, ootx_payloads_0_244, 
        ootx_payloads_0_188, n11209, n11800, ootx_payloads_0_187, n11208, 
        n2312, n11662, n22284, ootx_payloads_0_49, n11070, n11799, 
        ootx_payloads_0_186, n11207, n2604, n22685, n1405_c, n22462, 
        n22283, n2898, n2799, n22741, n2605, n22684, n22253, n22282, 
        n2192, n22586, n22252, n22227, n1406_c, n22461, n22216, 
        n22217, n2606, n22683, n3089, n22805, n2193, n22585, n22251, 
        n22281, n22250, n11727, n22226, n11661, ootx_payloads_0_48, 
        n11069, n11798, n1407_c, n22460, n2993, n22773, n2194, 
        n22584, n2899, n2800, n22740, n2607, n22682, ootx_payloads_0_185, 
        n11206, n23989, n23990, n22280, n1408_c, n22459, n22279, 
        n2608, n22681, ootx_payloads_0_243, n2900, n2801, n22739, 
        n22249, n22278, n22248, n2195, n22583, n22225, n11797, 
        ootx_payloads_0_242, n3012, n3011, n3010, n22903, n3009, 
        n30_adj_1907, n2999, n3005, n3006, n42_c, n2996, n3000, 
        n3001, n40_adj_1908, n2994, n3003, n3004, n45_c, n3007, 
        n44_c, n2995, n2997, n2998, n43_adj_1909, n3002, n47_c, 
        n1409_c, n25184, n22458, n2609, n25178, n22680, ootx_payloads_0_184, 
        n11205, ootx_payloads_0_76, n11097, n22247, n2196, n22582, 
        n22277, n22246, n11660, n22224, ootx_payloads_0_47, n11068, 
        n22215, n24110, n23992, n1410_c, n22457, n63_c, n3116, 
        n22842, n4731, n9989, ootx_payloads_0_241, n2610, n22679, 
        n2197, n22581, ootx_payloads_0_240, n93, n20098, n109, n3008, 
        n49_c, n1411_c, n22456, n22580, n11796, n1412_c, n22455, 
        n3090, n22804, n22772, ootx_payloads_0_183, n11204, n2901, 
        n2802, n22738, n2611, n22678, n22579, n112, n119, n22578, 
        n1301_c, n1334_c, n22454, n11795, n2612, n22677, ootx_payloads_0_182, 
        n11203, n22577, n117, n11659, n1302_c, n22453, n3, n23993, 
        n23994, n23996, n22576, n1303_c, n22452, ootx_payloads_0_227, 
        n11248, ootx_payloads_0_46, n11067, n2902, n2803, n22737, 
        n11794, n61_c, n22841, n22575, n1304_c, n22451, n22574, 
        n1305_c, n22450, ootx_payloads_0_181, n11202, n115, n2588, 
        n2489, n22676, n11793, ootx_payloads_0_180, n11201, n22573, 
        n1306_c, n22449, n2589, n2490, n22675, n22572, n110_adj_1911, 
        n1307_c, n22448, n11688, n3091, n22803, ootx_payloads_0_75, 
        n11096, n22771, n2903, n2804, n22736, n11658, n22571, 
        ootx_payloads_0_45, n11066, n11792, ootx_payloads_0_179, n11200;
    wire [5:0]sensor_state_switch_counter;   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(32[9:36])
    
    wire n37_adj_1914, n11726, ootx_payloads_0_226, n11247, n23995, 
        n11791, ootx_payloads_0_178, n11199, n107, n59_c, n22840, 
        n1308_c, n22447, n2590, n2491, n22674, n291, n22900, n4_adj_1917, 
        n24114, n9029, n30_adj_1918, n22276, n2591, n2492, n22673, 
        n22770, n25185, n22570, n22275, n2904, n2805, n22735, 
        n1309_c, n25186, n22446, n22245, n22244, n2493, n22672, 
        n2905, n2806, n22734, n22223, n2494, n22671, n22569, n1310_c, 
        n22445, n34_adj_1919, n32_adj_1920, n33_adj_1921, n31_adj_1922, 
        n24674, n24679, n24680, n271, n19257, n22273, n22568, 
        n22243, n22222, n22242, n1311_adj_1923, n22444, n22567, 
        n2495, n22670, n22272, n2496, n22669, n22271, n1312_adj_1925, 
        n22443, n2906, n2807, n22733, n22769, n6849, n23997, n23967, 
        n6_adj_1926, n7036, n22949, n22878, n24_adj_1927, n22877, 
        n23970, n2280, n22241, n22270, n2497, n22668, n22221, 
        n1994, n22566, n22240, n23775, n1995, n22565, n22239, 
        n1202_adj_1928, n22442, n22269, n2907, n2808, n22732, n2498, 
        n22667, n22220, n22238, n3092, n22802, n1203_adj_1929, n22441, 
        n2499, n22666, n1996, n22564, n16_adj_1930, n22_adj_1931, 
        n20_adj_1932, n24_adj_1933, n9196, n6_adj_1934, n22857, n10_adj_1935, 
        n6_adj_1936, n22268, n2908, n2809, n25180, n22731, n22267, 
        n11790, n1204_adj_1938, n22440, n2500, n22665, n57_c, n22839, 
        n1997, n22563, ootx_payloads_0_177, n11198, n11657, n1998, 
        n22562, n1205_adj_1940, n22439, ootx_payloads_0_44, n11065, 
        n11789, ootx_payloads_0_176, n11197, n11788, ootx_payloads_0_175, 
        n11196, n20_adj_1943, n43_adj_1944, n75, n103, n11656, ootx_payloads_0_43, 
        n11064, n11787, ootx_payloads_0_174, n11195, n11725, n11655, 
        ootx_payloads_0_42, n11063, n101, n11654, ootx_payloads_0_41, 
        n11062, n41_adj_1946, n234, n233, n11707, n73, n134_adj_1948, 
        n11786, ootx_payloads_0_173, n11194, n37_adj_1949, n262, n261, 
        n11653, ootx_payloads_0_40, n11061, n99, n11724, n11785, 
        ootx_payloads_0_172, n11193, n11652, ootx_payloads_0_39, n10995, 
        n11784, ootx_payloads_0_171, n11192, n11651, ootx_payloads_0_38, 
        n11020, n95, n11650, ootx_payloads_0_37, n10981, n11649, 
        ootx_payloads_0_225, n2501, n22664, ootx_payloads_0_36, n11022, 
        ootx_payloads_0_224, n168, n59_adj_1950, n252, n167, n11648, 
        n53_c, n13_adj_1951, n30_adj_1952, n3211, n3210, n22885, 
        n25_adj_1953, n27_adj_1954, n48_c, n15_adj_1955, n33_adj_1956, 
        n29_adj_1957, n35_adj_1958, n46_c, n41_adj_1959, n47_adj_1960, 
        n43_adj_1961, n47_adj_1962, n49_adj_1963, n51_c, n11, n45_adj_1964, 
        n17_adj_1965, n37_adj_1966, n19_adj_1967, n45_adj_1968, n44_adj_1969, 
        n21_adj_1970, n3209, n43_adj_1971, n54_c, n31_adj_1972, n55_c, 
        n39_adj_1973, n23_adj_1974, n49_adj_1975, n3215, ootx_payloads_0_35, 
        n10980, ootx_payloads_0_223, n11723, n11783, ootx_payloads_0_170, 
        n11191, n11647, ootx_payloads_0_34, n10985, ootx_payloads_0_222, 
        ootx_payloads_0_221, ootx_payloads_0_220, ootx_payloads_0_219, 
        n6_adj_1977, n11646, n26307, n6_adj_1979;
    wire [4:0]n5328;
    
    wire n24120, n24806, n24145, ootx_payloads_0_217, n1206_adj_1980, 
        n22438, n1999, n22561, ootx_payloads_0_33, n11000, ootx_payloads_0_216, 
        n93_adj_2014, n11782, n2000, n22560, n22838, n2909, n2810, 
        n22730, n1207_adj_2015, n22437, n22768, ootx_payloads_0_215, 
        ootx_payloads_0_169, n11190, n11645, ootx_payloads_0_214, n3093, 
        n22801, ootx_payloads_0_32, n10990, n22767, n251, n11687, 
        ootx_payloads_0_213, n2502, n22663, n2910, n2811, n22729, 
        n1208_adj_2017, n22436, ootx_payloads_0_212, n166_adj_2018, 
        n2001, n22559, n165, ootx_payloads_0_211, n11644, ootx_payloads_0_74, 
        n11095, n2503, n22662, ootx_payloads_0_31, n11017, n2002, 
        n22558, n11643, ootx_payloads_0_30, n11013, ootx_payloads_0_210, 
        n11781, ootx_payloads_0_168, n11189, ootx_payloads_0_209, n1209_adj_2021, 
        n22435, n11642, ootx_payloads_0_29, n11019, n2003, n22557, 
        n1210_adj_2023, n22434, n22837, n11641, ootx_payloads_0_28, 
        n11009, n11640, ootx_payloads_0_207, ootx_payloads_0_206, ootx_payloads_0_27, 
        n10982, ootx_payloads_0_205, ootx_payloads_0_204, n11780, n11246, 
        n3094, n22800, ootx_payloads_0_167, n11188, n22836, n11639, 
        ootx_payloads_0_26, n10983, n11245, n87, n11638, ootx_payloads_0_25, 
        n10984, n11779, ootx_payloads_0_166, n11187, n19283, n11637, 
        n11244, ootx_payloads_0_24, n10987, n11722, n35_adj_2030, 
        n164, n163, n1211_adj_2031, n22433, n2004, n22556, n2504, 
        n22661, n25219, n25222, n11721, n11636, n22835, ootx_payloads_0_23, 
        n10988, n11778, ootx_payloads_0_165, n11186, n2005, n22555, 
        n226, n1212_adj_2033, n22432, n22834, n23969, n2006, n22554, 
        n225, n11243, n11635, n2911, n2812, n22728, n2505, n22660, 
        n22766, n22237, ootx_payloads_0_22, n10989, n3095, n22799, 
        n22431, n83_adj_2035, n2912, n11634, n3096, n22798, ootx_payloads_0_21, 
        n10991, n11777, ootx_payloads_0_164, n11185, n11686, n11633, 
        ootx_payloads_0_20, n10992, n11706, n11632, n2007, n22553, 
        n22430, n22266, ootx_payloads_0_19, n10993, ootx_payloads_0_73, 
        n11094, n132, n2506, n22659, n2008, n22552, n22429, n60_adj_2038, 
        n11_adj_2039, n260, n259, n11631, ootx_payloads_0_18, n10994, 
        n2507, n22658, n2009, n22551, n22428, n2010, n22550, n22427, 
        n11776, ootx_payloads_0_163, n11184, n2786, n22727, n22214, 
        n11630, n2508, n22657, n2011, n22549, n22219, ootx_payloads_0_17, 
        n10996, n22426, n22236, n11629, ootx_payloads_0_16, n10997, 
        n2012, n22548, n22425, n2509, n22656, n11736, n11775, 
        ootx_payloads_0_162, n11183, n22424, n2787, n22726, n22547, 
        n22235, n2510, n22655, n22423, n22265, n22546, n22833, 
        n3097, n22797, n36_adj_2041, n22765, n11676, n170_adj_2042, 
        n19251, n22422, n2511, n22654, n172, n112_adj_2043, ootx_payloads_0_63, 
        n11084, n22545, n22218, n22544, n114_adj_2044, n116, n22421, 
        n22234, n2788, n22725, n22764, n11733, n120, n57_adj_2045, 
        n250, n249, n122_adj_2046;
    wire [30:0]n129;
    
    wire n2512, n22653, n22543, n124, n128, n22420, n11820, n22542, 
        n22419, n130_adj_2047, n2789, n22724, n22541, n22264, n11242, 
        n22418, n22652, n77, n22540, n22417, n218, n58_adj_2048, 
        n2790, n22723, n220, n22651, n22650, n22539, n22416, n11241, 
        n22538, n22263, n22415, n11228, n22537, n22414, n22233, 
        n22763, n11675, n22649, ootx_payloads_0_161, ootx_payloads_0_160, 
        n22536, n22413, n256, ootx_payloads_0_159, n2791, n22722, 
        ootx_payloads_0_158, n11732, n22648, n258, n22535, ootx_payloads_0_157, 
        n22534, ootx_payloads_0_156, ootx_payloads_0_155, ootx_payloads_0_154, 
        n22412, n22411, ootx_payloads_0_153, ootx_payloads_0_152, n22533, 
        n22647, n24676, n40_adj_2049, ootx_payloads_0_151, n22532, 
        n22410, ootx_payloads_0_150, n22721, n22409, n161, ootx_payloads_0_149, 
        n22646, ootx_payloads_0_148, n22531, n24682, n119_adj_2050, 
        ootx_payloads_0_147, ootx_payloads_0_146, n22530, n22408, n193_adj_2051, 
        n4_adj_2052, n257, n11240, ootx_payloads_0_145, n283, n223, 
        n256_adj_2053, n22645, n22407, ootx_payloads_0_144, ootx_payloads_0_143, 
        n11685, n169, n171, n3098, n22796, n24004, ootx_payloads_0_142, 
        ootx_payloads_0_141, ootx_payloads_0_140, n6_adj_2054, n22762, 
        n7, n118_adj_2055, n22406, n5, ootx_payloads_0_72, n11093, 
        n22720, n22529, data_N_1765, ootx_payloads_0_139, n22644, 
        ootx_payloads_0_138, ootx_payloads_0_137, ootx_payloads_0_136, 
        ootx_payloads_0_135, n22528, n22405, n22527, ootx_payloads_0_134, 
        ootx_payloads_0_133, ootx_payloads_0_132, ootx_payloads_0_131, 
        n22643, ootx_payloads_0_130, n22526, ootx_payloads_0_129, n22404, 
        n22403, ootx_payloads_0_128, n22525, ootx_payloads_0_127, n217, 
        n22719, n219, ootx_payloads_0_126, n22642, ootx_payloads_0_125, 
        n22524, n22402, ootx_payloads_0_124, n22523, n22401, n22641, 
        n22522, n22400, n22521, n22399, n18844, n22761, n11731, 
        n22718, n22760, n22640, n22520, n22398, n22519, n2276, 
        n10_adj_2057, n11713, n22639, n22518, n3099, n22795, n22397, 
        n22396, n255, n22517, n1631_adj_2058, n25199, n63_adj_2059, 
        n22395, n22832, n11628, n22717, n22638, ootx_payloads_0_15, 
        n10998, n22516, n22394, n11830, n22515, n22393, n11774, 
        n11829, n22637, n11182, ootx_payloads_0_62, n11083, n11828, 
        n22514, n3100, n22794, n22392, n22759, n11827, n11773, 
        n11181, n22513, n11627, ootx_payloads_0_14, n10999, n11826, 
        n3101, n22793, n11825, n22831, n11824, n22391, n22758, 
        n11705, n11823, n22636, n22716, n11822, n22390, n22355, 
        n3102, n22792, n22512, n22356, n11772, n22830, n11180, 
        n22635, n11626, n22511, n22354, n11819, n22389, ootx_payloads_0_13, 
        n11001, n22715, n11818, n11771, n11179, n11817, n22634, 
        n22510, n22388, n22353, n22714, n11704, n11625, ootx_payloads_0_12, 
        n11002, n25194, n22633, n22829, n22757, n22352, n11770, 
        n11178, n11624, ootx_payloads_0_11, n11003, n22828, n11623, 
        ootx_payloads_0_10, n11004, n11769, n22509, ootx_payloads_0_71, 
        n11177, ootx_payloads_0_70, n11622, n22387, ootx_payloads_0_9, 
        n11005, ootx_payloads_0_69, n22713, n22827, ootx_payloads_0_68, 
        n22632, ootx_payloads_0_67, ootx_payloads_0_66, ootx_payloads_0_65, 
        n65_c, n22508, n22351, ootx_payloads_0_64, n11703, n11621, 
        ootx_payloads_0_8, n11006, n11768, n11176, ootx_payloads_0_61, 
        n11620, n22631, n11730, ootx_payloads_0_60, ootx_payloads_0_7, 
        n11008, n11712, n22507;
    wire [5:0]n100;
    
    wire n22386;
    wire [15:0]n577;
    
    wire n22319, n22385, n4501, n22630, n22712, n11227, n11619, 
        n22506, ootx_payloads_0_6, n11010, n11767, n11684, n22318, 
        n22384, n11175, n22756, n11702, n11618, ootx_payloads_0_5, 
        n11014, n11766, n11174, n11617, ootx_payloads_0_4, n11015, 
        n22505, n22317, n11701, n11765, n11173, n11616, n22383, 
        n2291, n22629, n3103, n22791, n11092, ootx_payloads_0_3, 
        n11018, n22504, n11615, n22711, ootx_payloads_0_2, n11021, 
        n2292, n22628, n22382, n11700, n11764, n11172, n11614, 
        n22316, n22503, ootx_payloads_0_1, n11059, n2293, n22627, 
        n22826, n11613, ootx_payloads_0_0, n11060, n11763, n11171, 
        n11699, n22502, n22315, n11720, n11698, n22381, n11_adj_2070, 
        n22755, n22710, n2294, n22626, n12_adj_2072, n22501, n22314, 
        n22380, n11697, n2295, n22625, n11729, n25197, n22500, 
        n22379, n22313, n11683, n22709, n8_adj_2075, n9, n9_adj_2077, 
        n11762, n2296, n22624, n22499, n22378, n11170, n11696, 
        n10_adj_2079, n22623, n11091, n22498, n22377, n11695, n22312, 
        n22708, n11761, n11169, n11226, n22497, n22622, n22376, 
        n22311, n11760, n11168, n22375, n20123, n22621, n22707, 
        n1598_adj_2086, n22496, n22310, n11682, n22374, n1599_adj_2087, 
        n22495, n22620, n11012, n22825, n22309, n22824, n3104, 
        n22790, n22373, n1600_adj_2090, n22494, n22619, n22823, 
        n26_adj_2092, n42_adj_2093, n40_adj_2094, n41_adj_2095, n39_adj_2096, 
        n22891, n11759, n11167, n11090, n11758, n11757, n11756, 
        n11755, n11754, n11753, n11752, n11751, n11750, n11749, 
        n11748, n11747, n11746, n11745, n11744, n11743, n11742, 
        n11741, n11740, n11739, n11738, n11737, n11719, n11718, 
        n11717, n11716, n11715, n11711, n11710, n11709, n11694, 
        n11693, n11681, n11680, n11679, n11678, n11677, n11674, 
        n11673, n11089, n11166, n36_adj_2133, n11040, n22822, n11035, 
        n11030, n11039, n3105_adj_2136, n22789, n11026, n11034, 
        n22754, n22753, n11031, n11025, n11033, n11032, n11024, 
        n11023, n11238, n11037, n11028, n11036, n22706, n11029, 
        n22618, n44_adj_2137, n48_adj_2138, n11038, n11027, n11088, 
        n22372, n12_adj_2139, n22868, n11011, n11165, n11164, n19263, 
        n16_adj_2143, n17_adj_2144, n11163, n11284, n16_adj_2146, 
        n11162, n17_adj_2147, n11283, n15_adj_2148, n14_adj_2149, 
        n23991, n1601_adj_2150, n22493, n22308, n11161, n11160, 
        n22821, n11087, n11086, n11085, n11082, n11081, n11282, 
        n24564, n11281, n11280, n11279, n11278, n11277, n11276, 
        n11275, n11274, n11273, n11272, n11271, n11270, n11269, 
        n11268, n11267, n11266, n11265, n11264, n11263, n11262, 
        n11261, n11237, n11236, n11235, n11234, n11233, n11232, 
        n11231, n11230, n11225, n22617, n35_adj_2153, n22371, n11058, 
        n11159, n1602_adj_2154, n22492, n22307, n3106_adj_2155, n22788, 
        n11158, n22705, n22616, n22873, n14_adj_2156, n22370, n9_adj_2157, 
        n3112_c, n3111_adj_2158, n3110_adj_2159, n22889, n22491, n22306, 
        n18_adj_2160, n22942, n3108_adj_2161, n3109_adj_2162, n38_adj_2163, 
        n11157, n45_adj_2164, n22615, n28_adj_2165, n22369, n26_adj_2166, 
        n11156, n27_adj_2167, n3107_adj_2168, n42_adj_2169, n25_adj_2170, 
        n22820, n22490, n11155, n32_adj_2171, n19_adj_2172, n11154, 
        n11153, n22305, n22704, n22752, n11152, n18_adj_2173, n44_adj_2174, 
        n11151, n50_adj_2175, n11150, n48_adj_2177, n22614, n49_adj_2179, 
        n11149, n12_adj_2180, n47_adj_2181, n22368, n22489, n22304, 
        n26_adj_2182, n36_adj_2183, n22819, n11148, n22894, n24_adj_2184, 
        n11147, n22613, n11057, n23_adj_2185, n40_adj_2186, n22367, 
        n22488, n38_adj_2187, n39_adj_2188, n37_adj_2189, n22303, 
        n30_adj_2190, n22703, n40_adj_2191, n22787, n22612, n11056, 
        n22892, n38_adj_2192, n25_adj_2193, n44_adj_2194, n22366, 
        n11055, n42_adj_2195, n22487, n22302, n22611, n11054, n43_adj_2196, 
        n11053, n22365, n41_adj_2197, n22486, n22301, n6_adj_2198, 
        n11052, n19448, n18_adj_2199, n22786, n22818, n22702, n11051, 
        n16_adj_2200, n11050, n20_adj_2201, n11049, n22610, n22751, 
        n11048, n11047, n11046, n11042, n22364, n22485, n13338, 
        n13346, n22609, n22300, n22785, n22363, n22484, n23999, 
        n22299, n11146, n22608, n22948, n16_adj_2205, n22817, n22362, 
        n19_adj_2206, n18_adj_2207, n22_adj_2208, n22483, n11145, 
        n6_adj_2209, n19307, n30_adj_2210, n34_adj_2211, n32_adj_2212, 
        n33_adj_2213, n31_adj_2215, n22298, n22361, n22482, n22784, 
        n22816, n22701, n22297, n22607, n22750, n22360, n22783, 
        n22700, n22606, n24_adj_2226, n34_adj_2227, n32_adj_2228, 
        n22895, n22359, n22296, n38_adj_2229, n36_adj_2230, n22481, 
        n37_adj_2231, n35_adj_2232, n22605, n14_adj_2233, n22872, 
        n12_adj_2234, n16_adj_2235, n22480, n22295, n22358, n22699, 
        n22604, n22815, n22479, n22357, n22294, n28_adj_2237, n22814, 
        n22603, n31_adj_2238, n22947, n22_adj_2239, n30_adj_2240, 
        n34_adj_2241, n21_adj_2242;
    
    SB_LUT4 i6935_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_3), .I3(ootx_shift_registers_1_4), 
            .O(n11045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6935_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_1540_17_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n22601), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_355_20_lut (.I0(GND_net), .I1(counter_from_last_rise[18]), 
            .I2(GND_net), .I3(n22292), .O(n6333[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20515_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25183));
    defparam i20515_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE i671__i1 (.Q(\ootx_payload_o[1][0] ), .C(clock_c), .E(n2283), 
            .D(n2[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_CARRY mod_155_add_1071_12 (.CI(n22477), .I0(n1503), .I1(n1532), 
            .CO(n22478));
    SB_LUT4 mod_155_add_1942_23_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n22748), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_23_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n22697), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1808_23 (.CI(n22697), .I0(n2592), .I1(n2621), 
            .CO(n22698));
    SB_CARRY mod_155_add_1540_17 (.CI(n22601), .I0(n2198), .I1(n2225), 
            .CO(n22602));
    SB_CARRY add_355_20 (.CI(n22292), .I0(counter_from_last_rise[18]), .I1(GND_net), 
            .CO(n22293));
    SB_LUT4 i20530_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25198));
    defparam i20530_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6933_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_1), .I3(ootx_shift_registers_1_2), 
            .O(n11043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6933_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_355_19_lut (.I0(GND_net), .I1(counter_from_last_rise[17]), 
            .I2(GND_net), .I3(n22291), .O(n6333[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6130_4_lut_4_lut (.I0(n1119), .I1(\lighthouse[0] ), .I2(crc32s_N_1751), 
            .I3(n10243), .O(n1));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(153[22:32])
    defparam i6130_4_lut_4_lut.LUT_INIT = 16'hfd30;
    SB_LUT4 i6548_4_lut_4_lut (.I0(n1119), .I1(\lighthouse[0] ), .I2(n22972), 
            .I3(n1087), .O(n1_adj_1));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(153[22:32])
    defparam i6548_4_lut_4_lut.LUT_INIT = 16'h1f0f;
    SB_LUT4 mod_155_add_1071_11_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n22476), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1942_23 (.CI(n22748), .I0(n2792), .I1(n2819), 
            .CO(n22749));
    SB_LUT4 i7742_3_lut_4_lut (.I0(n1000), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1194), .O(n11852));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7742_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_19_i1_3_lut (.I0(payload_lengths_0_1), .I1(payload_lengths_1_1), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[1] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_19_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1540_16_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n22600), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_22_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n22696), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1071_11 (.CI(n22476), .I0(n1504), .I1(n1532), 
            .CO(n22477));
    SB_CARRY add_355_19 (.CI(n22291), .I0(counter_from_last_rise[17]), .I1(GND_net), 
            .CO(n22292));
    SB_LUT4 mod_155_add_2143_3_lut (.I0(n2851[1]), .I1(n2851[1]), .I2(n25181), 
            .I3(n22812), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1808_22 (.CI(n22696), .I0(n2593), .I1(n2621), 
            .CO(n22697));
    SB_LUT4 i6931_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(data), .I3(ootx_shift_registers_1_0), .O(n11041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6931_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY mod_155_add_1540_16 (.CI(n22600), .I0(n2199), .I1(n2225), 
            .CO(n22601));
    SB_LUT4 mod_155_add_1071_10_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n22475), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1540_15_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n22599), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1071_10 (.CI(n22475), .I0(n1505), .I1(n1532), 
            .CO(n22476));
    SB_LUT4 add_154_20_lut (.I0(GND_net), .I1(n2849[18]), .I2(GND_net), 
            .I3(n22261), .O(n2851[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2009_30_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n22782), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_30_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7150_3_lut_4_lut (.I0(n1000), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_239), .O(n11260));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7150_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_154_20 (.CI(n22261), .I0(n2849[18]), .I1(GND_net), .CO(n22262));
    SB_LUT4 mod_155_add_1942_22_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n22747), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_21_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n22695), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1540_15 (.CI(n22599), .I0(n2200), .I1(n2225), 
            .CO(n22600));
    SB_LUT4 Mux_29_i1_3_lut (.I0(bit_counters_0_7), .I1(bit_counters_1_7), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[7]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2143_3 (.CI(n22812), .I0(n2851[1]), .I1(n25181), 
            .CO(n22813));
    SB_LUT4 i6934_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_2), .I3(ootx_shift_registers_1_3), 
            .O(n11044));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6934_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 Mux_28_i1_3_lut (.I0(bit_counters_0_8), .I1(bit_counters_1_8), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[8]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_28_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1071_9_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n22474), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i647_648 (.Q(ootx_payloads_0_123), .C(clock_c), .D(n11144));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_27_i1_3_lut (.I0(bit_counters_0_9), .I1(bit_counters_1_9), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[9]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_27_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_3_lut (.I0(n2093), .I1(n2099), .I2(n2103), .I3(GND_net), 
            .O(n26));
    defparam i9_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut (.I0(n2098), .I1(n2104), .I2(n2097), .I3(n2105), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1540_14_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n22598), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_355_18_lut (.I0(GND_net), .I1(counter_from_last_rise[16]), 
            .I2(GND_net), .I3(n22290), .O(n6333[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(n2851[11]), .I1(n2112), .I2(n2111), .I3(n2110), 
            .O(n22941));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1071_9 (.CI(n22474), .I0(n1506), .I1(n1532), 
            .CO(n22475));
    SB_DFF i644_645 (.Q(ootx_payloads_0_122), .C(clock_c), .D(n11143));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i3_2_lut (.I0(n2096), .I1(n2102), .I2(GND_net), .I3(GND_net), 
            .O(n20_c));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 Mux_18_i1_3_lut (.I0(payload_lengths_0_2), .I1(payload_lengths_1_2), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[2] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_18_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut (.I0(n2100), .I1(n2101), .I2(n2108), .I3(n2107), 
            .O(n28_c));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n29), .I1(n2095), .I2(n26), .I3(n2106), .O(n32));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF i641_642 (.Q(ootx_payloads_0_121), .C(clock_c), .D(n11142));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_2009_29_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n22781), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut (.I0(ootx_payloads_N_1699[0]), .I1(n8941), .I2(n88), 
            .I3(GND_net), .O(n17_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(ootx_payloads_N_1699[0]), .I1(n8941), 
            .I2(n24018), .I3(\ootx_payloads_N_1699[4] ), .O(n13221));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff8;
    SB_DFF i638_639 (.Q(ootx_payloads_0_120), .C(clock_c), .D(n11141));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_adj_38 (.I0(reset_c), .I1(new_data), .I2(ootx_payloads_N_1744[0]), 
            .I3(GND_net), .O(n20112));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i1_2_lut_3_lut_adj_38.LUT_INIT = 16'hbfbf;
    SB_DFF i635_636 (.Q(ootx_payloads_0_119), .C(clock_c), .D(n11140));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1808_21 (.CI(n22695), .I0(n2594), .I1(n2621), 
            .CO(n22696));
    SB_LUT4 i3_4_lut_adj_39 (.I0(n2851[15]), .I1(n1712), .I2(n1711), .I3(n1710), 
            .O(n22946));
    defparam i3_4_lut_adj_39.LUT_INIT = 16'hfffe;
    SB_DFF i632_633 (.Q(ootx_payloads_0_118), .C(clock_c), .D(n11139));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i3_2_lut_adj_40 (.I0(n1699), .I1(n1706_adj_1810), .I2(GND_net), 
            .I3(GND_net), .O(n16));
    defparam i3_2_lut_adj_40.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(n22941), .I1(n2094), .I2(n2109), .I3(GND_net), 
            .O(n19_c));
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i9_4_lut (.I0(n1704), .I1(n1707), .I2(n1700), .I3(n1701), 
            .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF i629_630 (.Q(ootx_payloads_0_117), .C(clock_c), .D(n11138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i16_4_lut (.I0(n19_c), .I1(n32), .I2(n28_c), .I3(n20_c), 
            .O(n2126));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n22946), .I1(n1705), .I2(n1709), .I3(n1702), 
            .O(n20_adj_1811));
    defparam i7_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i11_4_lut_adj_41 (.I0(n1697), .I1(n22), .I2(n16), .I3(n1708), 
            .O(n24));
    defparam i11_4_lut_adj_41.LUT_INIT = 16'hfffe;
    SB_LUT4 Mux_26_i1_3_lut (.I0(bit_counters_0_10), .I1(bit_counters_1_10), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[10]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_26_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i626_627 (.Q(ootx_payloads_0_116), .C(clock_c), .D(n11137));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_adj_42 (.I0(reset_c), .I1(new_data), .I2(ootx_payloads_N_1744[1]), 
            .I3(GND_net), .O(n20105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i1_2_lut_3_lut_adj_42.LUT_INIT = 16'h4040;
    SB_CARRY mod_155_add_1540_14 (.CI(n22598), .I0(n2201), .I1(n2225), 
            .CO(n22599));
    SB_DFF i623_624 (.Q(ootx_payloads_0_115), .C(clock_c), .D(n11136));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_3_lut_4_lut (.I0(ootx_payloads_N_1744[1]), .I1(ootx_payloads_N_1744[0]), 
            .I2(n13221), .I3(data), .O(n23985));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[21:31])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i12_4_lut_adj_43 (.I0(n1698), .I1(n24), .I2(n20_adj_1811), 
            .I3(n1703), .O(n1730));
    defparam i12_4_lut_adj_43.LUT_INIT = 16'hfffe;
    SB_DFF i620_621 (.Q(ootx_payloads_0_114), .C(clock_c), .D(n11135));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i617_618 (.Q(ootx_payloads_0_113), .C(clock_c), .D(n11134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1071_8_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n22473), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_19_lut (.I0(GND_net), .I1(n2849[17]), .I2(GND_net), 
            .I3(n22260), .O(n2851[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20524_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25192));
    defparam i20524_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i614_615 (.Q(ootx_payloads_0_112), .C(clock_c), .D(n11133));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i611_612 (.Q(ootx_payloads_0_111), .C(clock_c), .D(n11132));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_17_i1_3_lut (.I0(payload_lengths_0_3), .I1(payload_lengths_1_3), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[3] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i608_609 (.Q(ootx_payloads_0_110), .C(clock_c), .D(n11131));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i605_606 (.Q(ootx_payloads_0_109), .C(clock_c), .D(n11130));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1540_13_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n22597), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_20_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[18]), 
            .I2(GND_net), .I3(n22231), .O(n337[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_44 (.I0(ootx_payloads_N_1744[1]), .I1(ootx_payloads_N_1744[0]), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n4));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[21:31])
    defparam i1_2_lut_3_lut_adj_44.LUT_INIT = 16'hb0b0;
    SB_DFF i602_603 (.Q(ootx_payloads_0_108), .C(clock_c), .D(n11129));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i2_3_lut_4_lut (.I0(\ootx_payloads_N_1699[4] ), .I1(n24018), 
            .I2(ootx_payloads_N_1744[1]), .I3(n20112), .O(n88));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF i599_600 (.Q(ootx_payloads_0_107), .C(clock_c), .D(n11128));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFR lighthouse_counter_639__i0 (.Q(\lighthouse[0] ), .C(clock_c), 
            .D(n69[0]), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    SB_DFF i596_597 (.Q(ootx_payloads_0_106), .C(clock_c), .D(n11127));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2009_29 (.CI(n22781), .I0(n2886), .I1(n2918), 
            .CO(n22782));
    SB_CARRY mod_155_add_1071_8 (.CI(n22473), .I0(n1507), .I1(n1532), 
            .CO(n22474));
    SB_LUT4 mod_155_add_2009_28_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n22780), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_28_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i593_594 (.Q(ootx_payloads_0_105), .C(clock_c), .D(n11126));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY add_66_20 (.CI(n22231), .I0(ootx_payloads_N_1699[18]), .I1(GND_net), 
            .CO(n22232));
    SB_LUT4 i7741_3_lut_4_lut (.I0(n998), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1195), .O(n11851));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7741_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_154_19 (.CI(n22260), .I0(n2849[17]), .I1(GND_net), .CO(n22261));
    SB_LUT4 i7149_3_lut_4_lut (.I0(n998), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_238), .O(n11259));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7149_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1942_22 (.CI(n22747), .I0(n2793), .I1(n2819), 
            .CO(n22748));
    SB_DFF i590_591 (.Q(ootx_payloads_0_104), .C(clock_c), .D(n11125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7740_3_lut_4_lut (.I0(n996), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1196), .O(n11850));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7740_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1808_20_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n22694), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1808_20 (.CI(n22694), .I0(n2595), .I1(n2621), 
            .CO(n22695));
    SB_LUT4 i20514_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25182));
    defparam i20514_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7148_3_lut_4_lut (.I0(n996), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_237), .O(n11258));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7148_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1540_13 (.CI(n22597), .I0(n2202), .I1(n2225), 
            .CO(n22598));
    SB_CARRY add_355_18 (.CI(n22290), .I0(counter_from_last_rise[16]), .I1(GND_net), 
            .CO(n22291));
    SB_LUT4 mod_155_add_1071_7_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n22472), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_18_lut (.I0(GND_net), .I1(n2849[16]), .I2(GND_net), 
            .I3(n22259), .O(n2851[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7739_3_lut_4_lut (.I0(n994), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1197), .O(n11849));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7739_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1540_12_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n22596), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1071_7 (.CI(n22472), .I0(n1508), .I1(n1532), 
            .CO(n22473));
    SB_CARRY mod_155_add_2143_2 (.CI(VCC_net), .I0(n2851[0]), .I1(VCC_net), 
            .CO(n22812));
    SB_CARRY mod_155_add_2009_28 (.CI(n22780), .I0(n2887), .I1(n2918), 
            .CO(n22781));
    SB_LUT4 mod_155_add_1808_19_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n22693), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_18 (.CI(n22259), .I0(n2849[16]), .I1(GND_net), .CO(n22260));
    SB_CARRY mod_155_add_1540_12 (.CI(n22596), .I0(n2203), .I1(n2225), 
            .CO(n22597));
    SB_LUT4 mod_155_add_1071_6_lut (.I0(n1509), .I1(n1509), .I2(n25177), 
            .I3(n22471), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_355_17_lut (.I0(GND_net), .I1(counter_from_last_rise[15]), 
            .I2(GND_net), .I3(n22289), .O(n6333[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7147_3_lut_4_lut (.I0(n994), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_236), .O(n11257));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7147_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1540_11_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n22595), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_17_lut (.I0(GND_net), .I1(n2849[15]), .I2(GND_net), 
            .I3(n22258), .O(n2851[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1071_6 (.CI(n22471), .I0(n1509), .I1(n25177), 
            .CO(n22472));
    SB_LUT4 i7738_3_lut_4_lut (.I0(n992), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1198), .O(n11848));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7738_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_66_19_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[17]), 
            .I2(GND_net), .I3(n22230), .O(n337[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2009_27_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n22779), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2076_31_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n22811), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_31_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2009_27 (.CI(n22779), .I0(n2888), .I1(n2918), 
            .CO(n22780));
    SB_LUT4 i7146_3_lut_4_lut (.I0(n992), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_235), .O(n11256));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7146_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1942_21_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n22746), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_19 (.CI(n22230), .I0(ootx_payloads_N_1699[17]), .I1(GND_net), 
            .CO(n22231));
    SB_CARRY add_154_17 (.CI(n22258), .I0(n2849[15]), .I1(GND_net), .CO(n22259));
    SB_LUT4 i7033_3_lut_4_lut (.I0(n766), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_122), .O(n11143));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7033_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1808_19 (.CI(n22693), .I0(n2596), .I1(n2621), 
            .CO(n22694));
    SB_CARRY mod_155_add_1540_11 (.CI(n22595), .I0(n2204), .I1(n2225), 
            .CO(n22596));
    SB_LUT4 mod_155_add_2009_26_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n22778), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7625_3_lut_4_lut (.I0(n766), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1311), .O(n11735));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7625_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_45 (.I0(n13), .I1(n24018), .I2(n9498), 
            .I3(n118), .O(crc32s_N_1751));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam i2_3_lut_4_lut_adj_45.LUT_INIT = 16'h1000;
    SB_LUT4 i7737_3_lut_4_lut (.I0(n990), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1199), .O(n11847));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7737_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1942_21 (.CI(n22746), .I0(n2794), .I1(n2819), 
            .CO(n22747));
    SB_LUT4 mod_155_add_1071_5_lut (.I0(n1510), .I1(n1510), .I2(n1532), 
            .I3(n22470), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7145_3_lut_4_lut (.I0(n990), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_234), .O(n11255));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7145_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1540_10_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n22594), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_18_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n22692), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1071_5 (.CI(n22470), .I0(n1510), .I1(n1532), 
            .CO(n22471));
    SB_LUT4 i20528_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25196));
    defparam i20528_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_155_add_1808_18 (.CI(n22692), .I0(n2597), .I1(n2621), 
            .CO(n22693));
    SB_LUT4 i9429_3_lut (.I0(n2851[24]), .I1(n71[24]), .I2(n839), .I3(GND_net), 
            .O(n912_c));
    defparam i9429_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1540_10 (.CI(n22594), .I0(n2205), .I1(n2225), 
            .CO(n22595));
    SB_CARRY add_355_17 (.CI(n22289), .I0(counter_from_last_rise[15]), .I1(GND_net), 
            .CO(n22290));
    SB_LUT4 i3_4_lut_adj_46 (.I0(n2851[14]), .I1(n1812), .I2(n1811), .I3(n1810), 
            .O(n22945));
    defparam i3_4_lut_adj_46.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1071_4_lut (.I0(n1511), .I1(n1511), .I2(n1532), 
            .I3(n22469), .O(n1610)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_355_16_lut (.I0(GND_net), .I1(counter_from_last_rise[14]), 
            .I2(GND_net), .I3(n22288), .O(n6333[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1540_9_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n22593), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_17_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n22691), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7736_3_lut_4_lut (.I0(n988), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1200), .O(n11846));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7736_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1071_4 (.CI(n22469), .I0(n1511), .I1(n1532), 
            .CO(n22470));
    SB_LUT4 i4_3_lut (.I0(n1799), .I1(n22945), .I2(n1809), .I3(GND_net), 
            .O(n18));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i7144_3_lut_4_lut (.I0(n988), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_233), .O(n11254));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7144_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut (.I0(n1805), .I1(n1802), .I2(n1803), .I3(n1797), 
            .O(n24_adj_1812));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1807), .I1(n1796), .I2(n1806), .I3(n1800), 
            .O(n22_adj_1813));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1942_20_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n22745), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_16 (.CI(n22288), .I0(counter_from_last_rise[14]), .I1(GND_net), 
            .CO(n22289));
    SB_LUT4 i6672_4_lut_4_lut (.I0(n1119), .I1(\lighthouse[0] ), .I2(n72[1]), 
            .I3(n1087), .O(n1_adj_2));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(153[22:32])
    defparam i6672_4_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_CARRY mod_155_add_1808_17 (.CI(n22691), .I0(n2598), .I1(n2621), 
            .CO(n22692));
    SB_LUT4 i12_4_lut_adj_47 (.I0(n1808), .I1(n24_adj_1812), .I2(n18), 
            .I3(n1801), .O(n26_adj_1815));
    defparam i12_4_lut_adj_47.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n1804), .I1(n26_adj_1815), .I2(n22_adj_1813), 
            .I3(n1798), .O(n1829));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1540_9 (.CI(n22593), .I0(n2206), .I1(n2225), 
            .CO(n22594));
    SB_LUT4 add_355_15_lut (.I0(GND_net), .I1(counter_from_last_rise[13]), 
            .I2(GND_net), .I3(n22287), .O(n6333[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1071_3_lut (.I0(n1512), .I1(n1512), .I2(n1532), 
            .I3(n22468), .O(n1611)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_3_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1942_20 (.CI(n22745), .I0(n2795), .I1(n2819), 
            .CO(n22746));
    SB_LUT4 i3_4_lut_4_lut (.I0(n1119), .I1(\lighthouse[0] ), .I2(n72[1]), 
            .I3(n24028), .O(n9797));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(153[22:32])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 i20462_2_lut (.I0(n23974), .I1(data), .I2(GND_net), .I3(GND_net), 
            .O(n24829));
    defparam i20462_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i587_588 (.Q(ootx_payloads_0_103), .C(clock_c), .D(n11124));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_2076_30_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n22810), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_30_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1540_8_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n22592), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i584_585 (.Q(ootx_payloads_0_102), .C(clock_c), .D(n11123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i9426_3_lut (.I0(n811), .I1(n71[26]), .I2(n839), .I3(GND_net), 
            .O(n910_c));
    defparam i9426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20527_1_lut (.I0(n938_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25195));
    defparam i20527_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i581_582 (.Q(ootx_payloads_0_101), .C(clock_c), .D(n11122));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i578_579 (.Q(ootx_payloads_0_100), .C(clock_c), .D(n11121));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2009_26 (.CI(n22778), .I0(n2889), .I1(n2918), 
            .CO(n22779));
    SB_DFF i575_576 (.Q(ootx_payloads_0_99), .C(clock_c), .D(n11120));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1071_3 (.CI(n22468), .I0(n1512), .I1(n1532), 
            .CO(n22469));
    SB_DFFE counter_from_last_rise__i0 (.Q(counter_from_last_rise[0]), .C(clock_c), 
            .E(VCC_net), .D(n8));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 mod_155_add_1808_16_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n22690), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_17_i1_3_lut_adj_48 (.I0(bit_counters_0_19), .I1(bit_counters_1_19), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[19]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_17_i1_3_lut_adj_48.LUT_INIT = 16'hcaca;
    SB_DFFE data_counters_0_0_c (.Q(data_counters_0_0), .C(clock_c), .E(VCC_net), 
            .D(n23003));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_1_c (.Q(data_counters_0_1), .C(clock_c), .E(VCC_net), 
            .D(n23005));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_2_c (.Q(data_counters_0_2), .C(clock_c), .E(VCC_net), 
            .D(n23007));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_3_c (.Q(data_counters_0_3), .C(clock_c), .E(VCC_net), 
            .D(n23009));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_4_c (.Q(data_counters_0_4), .C(clock_c), .E(VCC_net), 
            .D(n23011));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_5_c (.Q(data_counters_0_5), .C(clock_c), .E(VCC_net), 
            .D(n23013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_6_c (.Q(data_counters_0_6), .C(clock_c), .E(VCC_net), 
            .D(n23015));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_7_c (.Q(data_counters_0_7), .C(clock_c), .E(VCC_net), 
            .D(n23017));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_8_c (.Q(data_counters_0_8), .C(clock_c), .E(VCC_net), 
            .D(n23019));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_9_c (.Q(data_counters_0_9), .C(clock_c), .E(VCC_net), 
            .D(n23021));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_10_c (.Q(data_counters_0_10), .C(clock_c), .E(VCC_net), 
            .D(n23023));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_LUT4 i6244_4_lut_4_lut (.I0(n1119), .I1(\lighthouse[0] ), .I2(crc32s_N_1751), 
            .I3(n10357), .O(n1_adj_3));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(153[22:32])
    defparam i6244_4_lut_4_lut.LUT_INIT = 16'hf7c0;
    SB_DFFE data_counters_0_11_c (.Q(data_counters_0_11), .C(clock_c), .E(VCC_net), 
            .D(n23025));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_12_c (.Q(data_counters_0_12), .C(clock_c), .E(VCC_net), 
            .D(n23027));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_13_c (.Q(data_counters_0_13), .C(clock_c), .E(VCC_net), 
            .D(n23029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_14_c (.Q(data_counters_0_14), .C(clock_c), .E(VCC_net), 
            .D(n23031));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_15_c (.Q(data_counters_0_15), .C(clock_c), .E(VCC_net), 
            .D(n23033));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_16_c (.Q(data_counters_0_16), .C(clock_c), .E(VCC_net), 
            .D(n23035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_17_c (.Q(data_counters_0_17), .C(clock_c), .E(VCC_net), 
            .D(n23037));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_18_c (.Q(data_counters_0_18), .C(clock_c), .E(VCC_net), 
            .D(n23039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_19_c (.Q(data_counters_0_19), .C(clock_c), .E(VCC_net), 
            .D(n23041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_20_c (.Q(data_counters_0_20), .C(clock_c), .E(VCC_net), 
            .D(n23043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_21_c (.Q(data_counters_0_21), .C(clock_c), .E(VCC_net), 
            .D(n23045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_22_c (.Q(data_counters_0_22), .C(clock_c), .E(VCC_net), 
            .D(n23047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_23_c (.Q(data_counters_0_23), .C(clock_c), .E(VCC_net), 
            .D(n23049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_24_c (.Q(data_counters_0_24), .C(clock_c), .E(VCC_net), 
            .D(n23051));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_25_c (.Q(data_counters_0_25), .C(clock_c), .E(VCC_net), 
            .D(n23053));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_26_c (.Q(data_counters_0_26), .C(clock_c), .E(VCC_net), 
            .D(n23055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_27_c (.Q(data_counters_0_27), .C(clock_c), .E(VCC_net), 
            .D(n23057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_28_c (.Q(data_counters_0_28), .C(clock_c), .E(VCC_net), 
            .D(n23059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_29_c (.Q(data_counters_0_29), .C(clock_c), .E(VCC_net), 
            .D(n23061));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_0_30_c (.Q(data_counters_0_30), .C(clock_c), .E(VCC_net), 
            .D(n23063));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_0_c (.Q(data_counters_1_0), .C(clock_c), .E(VCC_net), 
            .D(n23065));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_1_c (.Q(data_counters_1_1), .C(clock_c), .E(VCC_net), 
            .D(n23067));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_2_c (.Q(data_counters_1_2), .C(clock_c), .E(VCC_net), 
            .D(n23069));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_3_c (.Q(data_counters_1_3), .C(clock_c), .E(VCC_net), 
            .D(n23071));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_4_c (.Q(data_counters_1_4), .C(clock_c), .E(VCC_net), 
            .D(n23073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_5_c (.Q(data_counters_1_5), .C(clock_c), .E(VCC_net), 
            .D(n23075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_6_c (.Q(data_counters_1_6), .C(clock_c), .E(VCC_net), 
            .D(n23077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_7_c (.Q(data_counters_1_7), .C(clock_c), .E(VCC_net), 
            .D(n23079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_8_c (.Q(data_counters_1_8), .C(clock_c), .E(VCC_net), 
            .D(n23081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_9_c (.Q(data_counters_1_9), .C(clock_c), .E(VCC_net), 
            .D(n23083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_10_c (.Q(data_counters_1_10), .C(clock_c), .E(VCC_net), 
            .D(n23085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_11_c (.Q(data_counters_1_11), .C(clock_c), .E(VCC_net), 
            .D(n23087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_12_c (.Q(data_counters_1_12), .C(clock_c), .E(VCC_net), 
            .D(n23089));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_13_c (.Q(data_counters_1_13), .C(clock_c), .E(VCC_net), 
            .D(n23091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_14_c (.Q(data_counters_1_14), .C(clock_c), .E(VCC_net), 
            .D(n23093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_15_c (.Q(data_counters_1_15), .C(clock_c), .E(VCC_net), 
            .D(n23095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_16_c (.Q(data_counters_1_16), .C(clock_c), .E(VCC_net), 
            .D(n23097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_17_c (.Q(data_counters_1_17), .C(clock_c), .E(VCC_net), 
            .D(n23099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_18_c (.Q(data_counters_1_18), .C(clock_c), .E(VCC_net), 
            .D(n23101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_19_c (.Q(data_counters_1_19), .C(clock_c), .E(VCC_net), 
            .D(n23103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_20_c (.Q(data_counters_1_20), .C(clock_c), .E(VCC_net), 
            .D(n23105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_21_c (.Q(data_counters_1_21), .C(clock_c), .E(VCC_net), 
            .D(n23107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_22_c (.Q(data_counters_1_22), .C(clock_c), .E(VCC_net), 
            .D(n23109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_23_c (.Q(data_counters_1_23), .C(clock_c), .E(VCC_net), 
            .D(n23111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_24_c (.Q(data_counters_1_24), .C(clock_c), .E(VCC_net), 
            .D(n23113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_25_c (.Q(data_counters_1_25), .C(clock_c), .E(VCC_net), 
            .D(n23115));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_26_c (.Q(data_counters_1_26), .C(clock_c), .E(VCC_net), 
            .D(n23117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_27_c (.Q(data_counters_1_27), .C(clock_c), .E(VCC_net), 
            .D(n23119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_28_c (.Q(data_counters_1_28), .C(clock_c), .E(VCC_net), 
            .D(n23121));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_29_c (.Q(data_counters_1_29), .C(clock_c), .E(VCC_net), 
            .D(n23123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE data_counters_1_30_c (.Q(data_counters_1_30), .C(clock_c), .E(VCC_net), 
            .D(n23125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    SB_DFFE bit_counters_0_0_c (.Q(bit_counters_0_0), .C(clock_c), .E(VCC_net), 
            .D(n23475));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_1_c (.Q(bit_counters_0_1), .C(clock_c), .E(VCC_net), 
            .D(n23477));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_2_c (.Q(bit_counters_0_2), .C(clock_c), .E(VCC_net), 
            .D(n23479));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_3_c (.Q(bit_counters_0_3), .C(clock_c), .E(VCC_net), 
            .D(n23481));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_4_c (.Q(bit_counters_0_4), .C(clock_c), .E(VCC_net), 
            .D(n23483));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_5_c (.Q(bit_counters_0_5), .C(clock_c), .E(VCC_net), 
            .D(n23485));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_6_c (.Q(bit_counters_0_6), .C(clock_c), .E(VCC_net), 
            .D(n23487));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_7_c (.Q(bit_counters_0_7), .C(clock_c), .E(VCC_net), 
            .D(n23489));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_8_c (.Q(bit_counters_0_8), .C(clock_c), .E(VCC_net), 
            .D(n23491));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_9_c (.Q(bit_counters_0_9), .C(clock_c), .E(VCC_net), 
            .D(n23493));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_10_c (.Q(bit_counters_0_10), .C(clock_c), .E(VCC_net), 
            .D(n23495));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_11_c (.Q(bit_counters_0_11), .C(clock_c), .E(VCC_net), 
            .D(n23497));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_12_c (.Q(bit_counters_0_12), .C(clock_c), .E(VCC_net), 
            .D(n23499));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_13_c (.Q(bit_counters_0_13), .C(clock_c), .E(VCC_net), 
            .D(n23501));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_14_c (.Q(bit_counters_0_14), .C(clock_c), .E(VCC_net), 
            .D(n23503));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_15_c (.Q(bit_counters_0_15), .C(clock_c), .E(VCC_net), 
            .D(n23505));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_16_c (.Q(bit_counters_0_16), .C(clock_c), .E(VCC_net), 
            .D(n23507));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_17_c (.Q(bit_counters_0_17), .C(clock_c), .E(VCC_net), 
            .D(n23509));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_18_c (.Q(bit_counters_0_18), .C(clock_c), .E(VCC_net), 
            .D(n23469));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_19_c (.Q(bit_counters_0_19), .C(clock_c), .E(VCC_net), 
            .D(n23463));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_20_c (.Q(bit_counters_0_20), .C(clock_c), .E(VCC_net), 
            .D(n23457));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_21_c (.Q(bit_counters_0_21), .C(clock_c), .E(VCC_net), 
            .D(n23451));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_22_c (.Q(bit_counters_0_22), .C(clock_c), .E(VCC_net), 
            .D(n23445));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_23_c (.Q(bit_counters_0_23), .C(clock_c), .E(VCC_net), 
            .D(n23439));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_24_c (.Q(bit_counters_0_24), .C(clock_c), .E(VCC_net), 
            .D(n23433));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_25_c (.Q(bit_counters_0_25), .C(clock_c), .E(VCC_net), 
            .D(n23427));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_26_c (.Q(bit_counters_0_26), .C(clock_c), .E(VCC_net), 
            .D(n23421));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_27_c (.Q(bit_counters_0_27), .C(clock_c), .E(VCC_net), 
            .D(n23415));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_28_c (.Q(bit_counters_0_28), .C(clock_c), .E(VCC_net), 
            .D(n23409));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_29_c (.Q(bit_counters_0_29), .C(clock_c), .E(VCC_net), 
            .D(n23399));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_0_30_c (.Q(bit_counters_0_30), .C(clock_c), .E(VCC_net), 
            .D(n23389));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_0_c (.Q(bit_counters_1_0), .C(clock_c), .E(VCC_net), 
            .D(n23511));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_1_c (.Q(bit_counters_1_1), .C(clock_c), .E(VCC_net), 
            .D(n23513));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_2_c (.Q(bit_counters_1_2), .C(clock_c), .E(VCC_net), 
            .D(n23515));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_3_c (.Q(bit_counters_1_3), .C(clock_c), .E(VCC_net), 
            .D(n23517));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_4_c (.Q(bit_counters_1_4), .C(clock_c), .E(VCC_net), 
            .D(n23519));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_5_c (.Q(bit_counters_1_5), .C(clock_c), .E(VCC_net), 
            .D(n23521));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_6_c (.Q(bit_counters_1_6), .C(clock_c), .E(VCC_net), 
            .D(n23523));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_7_c (.Q(bit_counters_1_7), .C(clock_c), .E(VCC_net), 
            .D(n23525));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_8_c (.Q(bit_counters_1_8), .C(clock_c), .E(VCC_net), 
            .D(n23527));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_9_c (.Q(bit_counters_1_9), .C(clock_c), .E(VCC_net), 
            .D(n23529));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_10_c (.Q(bit_counters_1_10), .C(clock_c), .E(VCC_net), 
            .D(n23531));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_11_c (.Q(bit_counters_1_11), .C(clock_c), .E(VCC_net), 
            .D(n23533));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_12_c (.Q(bit_counters_1_12), .C(clock_c), .E(VCC_net), 
            .D(n23535));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_13_c (.Q(bit_counters_1_13), .C(clock_c), .E(VCC_net), 
            .D(n23537));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_14_c (.Q(bit_counters_1_14), .C(clock_c), .E(VCC_net), 
            .D(n23539));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_15_c (.Q(bit_counters_1_15), .C(clock_c), .E(VCC_net), 
            .D(n23541));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_16_c (.Q(bit_counters_1_16), .C(clock_c), .E(VCC_net), 
            .D(n23543));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_17_c (.Q(bit_counters_1_17), .C(clock_c), .E(VCC_net), 
            .D(n23545));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_18_c (.Q(bit_counters_1_18), .C(clock_c), .E(VCC_net), 
            .D(n23471));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_19_c (.Q(bit_counters_1_19), .C(clock_c), .E(VCC_net), 
            .D(n23465));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_20_c (.Q(bit_counters_1_20), .C(clock_c), .E(VCC_net), 
            .D(n23459));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_21_c (.Q(bit_counters_1_21), .C(clock_c), .E(VCC_net), 
            .D(n23453));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_22_c (.Q(bit_counters_1_22), .C(clock_c), .E(VCC_net), 
            .D(n23447));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_23_c (.Q(bit_counters_1_23), .C(clock_c), .E(VCC_net), 
            .D(n23441));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_24_c (.Q(bit_counters_1_24), .C(clock_c), .E(VCC_net), 
            .D(n23435));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_25_c (.Q(bit_counters_1_25), .C(clock_c), .E(VCC_net), 
            .D(n23429));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_26_c (.Q(bit_counters_1_26), .C(clock_c), .E(VCC_net), 
            .D(n23423));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_27_c (.Q(bit_counters_1_27), .C(clock_c), .E(VCC_net), 
            .D(n23417));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_LUT4 i9428_3_lut (.I0(n809), .I1(n71[28]), .I2(n839), .I3(GND_net), 
            .O(n908_c));
    defparam i9428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9430_3_lut (.I0(n808_c), .I1(n71[29]), .I2(n839), .I3(GND_net), 
            .O(n907));
    defparam i9430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1942_19_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n22744), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1808_16 (.CI(n22690), .I0(n2599), .I1(n2621), 
            .CO(n22691));
    SB_CARRY add_355_15 (.CI(n22287), .I0(counter_from_last_rise[13]), .I1(GND_net), 
            .CO(n22288));
    SB_LUT4 i20523_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25191));
    defparam i20523_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_155_add_2076_30 (.CI(n22810), .I0(n2985), .I1(n3017), 
            .CO(n22811));
    SB_CARRY mod_155_add_1540_8 (.CI(n22592), .I0(n2207), .I1(n2225), 
            .CO(n22593));
    SB_LUT4 add_154_16_lut (.I0(GND_net), .I1(n2849[14]), .I2(GND_net), 
            .I3(n22257), .O(n2851[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9427_3_lut (.I0(n807), .I1(n71[30]), .I2(n839), .I3(GND_net), 
            .O(n906_c));
    defparam i9427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_i543_3_lut (.I0(n2851[25]), .I1(n773[25]), .I2(n740_c), 
            .I3(GND_net), .O(n812_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_i541_3_lut (.I0(n711), .I1(n773[27]), .I2(n740_c), 
            .I3(GND_net), .O(n810_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1071_2_lut (.I0(n2851[17]), .I1(n2851[17]), .I2(n25177), 
            .I3(VCC_net), .O(n1612)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_i608_3_lut (.I0(n810_c), .I1(n71[27]), .I2(n839), 
            .I3(GND_net), .O(n909));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_i610_3_lut (.I0(n812_c), .I1(n71[25]), .I2(n839), 
            .I3(GND_net), .O(n911));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7735_3_lut_4_lut (.I0(n986), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1201), .O(n11845));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7735_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_i539_3_lut (.I0(n709), .I1(n773[29]), .I2(n740_c), 
            .I3(GND_net), .O(n808_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_i538_3_lut (.I0(n708_c), .I1(n773[30]), .I2(n740_c), 
            .I3(GND_net), .O(n807));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7143_3_lut_4_lut (.I0(n986), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_232), .O(n11253));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7143_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i51_4_lut (.I0(\lighthouse[0] ), .I1(n24829), .I2(ootx_payloads_N_1744[0]), 
            .I3(n35), .O(n27));
    defparam i51_4_lut.LUT_INIT = 16'hc0c5;
    SB_DFFE bit_counters_1_28_c (.Q(bit_counters_1_28), .C(clock_c), .E(VCC_net), 
            .D(n23411));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_29_c (.Q(bit_counters_1_29), .C(clock_c), .E(VCC_net), 
            .D(n23401));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE bit_counters_1_30_c (.Q(bit_counters_1_30), .C(clock_c), .E(VCC_net), 
            .D(n23391));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(56[9:21])
    SB_DFFE new_data_477 (.Q(new_data), .C(clock_c), .E(VCC_net), .D(n23697));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE i24_25 (.Q(payload_lengths_0_0), .C(clock_c), .E(VCC_net), 
            .D(n23639));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i88_89 (.Q(payload_lengths_1_0), .C(clock_c), .E(VCC_net), 
            .D(n23641));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE counter_from_last_rise__i1 (.Q(counter_from_last_rise[1]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_4));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i2 (.Q(counter_from_last_rise[2]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_5));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 mod_155_i542_3_lut (.I0(n712_c), .I1(n773[26]), .I2(n740_c), 
            .I3(GND_net), .O(n811));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i542_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE counter_from_last_rise__i3 (.Q(counter_from_last_rise[3]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_6));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE i28_29 (.Q(payload_lengths_0_1), .C(clock_c), .E(n24097), 
            .D(n58_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_LUT4 mod_155_add_2076_29_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n22809), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_i472_3_lut (.I0(n610_c), .I1(n89[29]), .I2(n641), 
            .I3(GND_net), .O(n709));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i472_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE i32_33 (.Q(payload_lengths_0_2), .C(clock_c), .E(n24124), 
            .D(n62_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_LUT4 mod_155_add_1540_7_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n22591), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE i36_37 (.Q(payload_lengths_0_3), .C(clock_c), .E(n24095), 
            .D(n66_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i40_41 (.Q(payload_lengths_0_4), .C(clock_c), .E(n24093), 
            .D(n70));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i44_45 (.Q(payload_lengths_0_5), .C(clock_c), .E(n24091), 
            .D(n74));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFF i572_573 (.Q(ootx_payloads_0_98), .C(clock_c), .D(n11119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFE i48_49 (.Q(payload_lengths_0_6), .C(clock_c), .E(n24089), 
            .D(n78));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i52_53 (.Q(payload_lengths_0_7), .C(clock_c), .E(n24087), 
            .D(n82));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i56_57 (.Q(payload_lengths_0_8), .C(clock_c), .E(n24085), 
            .D(n86));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i60_61 (.Q(payload_lengths_0_9), .C(clock_c), .E(n24083), 
            .D(n90));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i64_65 (.Q(payload_lengths_0_10), .C(clock_c), .E(n24081), 
            .D(n94));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i68_69 (.Q(payload_lengths_0_11), .C(clock_c), .E(n24079), 
            .D(n98));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i72_73 (.Q(payload_lengths_0_12), .C(clock_c), .E(n24077), 
            .D(n102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i76_77 (.Q(payload_lengths_0_13), .C(clock_c), .E(n24075), 
            .D(n106));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFF i569_570 (.Q(ootx_payloads_0_97), .C(clock_c), .D(n11118));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFE i80_81 (.Q(payload_lengths_0_14), .C(clock_c), .E(n24073), 
            .D(n110));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i84_85 (.Q(payload_lengths_0_15), .C(clock_c), .E(n24071), 
            .D(n114));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i92_93 (.Q(payload_lengths_1_1), .C(clock_c), .E(n24069), 
            .D(n122));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_LUT4 mod_155_i471_3_lut (.I0(n609), .I1(n89[30]), .I2(n641), .I3(GND_net), 
            .O(n708_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i471_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE i96_97 (.Q(payload_lengths_1_2), .C(clock_c), .E(n24067), 
            .D(n126));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_LUT4 i1338_2_lut (.I0(n2851[29]), .I1(n58_adj_1820), .I2(GND_net), 
            .I3(GND_net), .O(n60_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i1338_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE i100_101 (.Q(payload_lengths_1_3), .C(clock_c), .E(n24065), 
            .D(n130));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i104_105 (.Q(payload_lengths_1_4), .C(clock_c), .E(n24063), 
            .D(n134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i108_109 (.Q(payload_lengths_1_5), .C(clock_c), .E(n24061), 
            .D(n138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFF i566_567 (.Q(ootx_payloads_0_96), .C(clock_c), .D(n11117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFE i112_113 (.Q(payload_lengths_1_6), .C(clock_c), .E(n24059), 
            .D(n142));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i116_117 (.Q(payload_lengths_1_7), .C(clock_c), .E(n24057), 
            .D(n146));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i120_121 (.Q(payload_lengths_1_8), .C(clock_c), .E(n24055), 
            .D(n150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i124_125 (.Q(payload_lengths_1_9), .C(clock_c), .E(n24053), 
            .D(n154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i128_129 (.Q(payload_lengths_1_10), .C(clock_c), .E(n24051), 
            .D(n158));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i132_133 (.Q(payload_lengths_1_11), .C(clock_c), .E(n24049), 
            .D(n162));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i136_137 (.Q(payload_lengths_1_12), .C(clock_c), .E(n24047), 
            .D(n166));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_CARRY mod_155_add_1071_2 (.CI(VCC_net), .I0(n2851[17]), .I1(n25177), 
            .CO(n22468));
    SB_DFFE i140_141 (.Q(payload_lengths_1_13), .C(clock_c), .E(n24045), 
            .D(n170));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFF i563_564 (.Q(ootx_payloads_0_95), .C(clock_c), .D(n11116));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFE counter_from_nskip_rise_640__i0 (.Q(counter_from_nskip_rise[0]), 
            .C(clock_c), .E(n2282), .D(n91[0]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE i144_145 (.Q(payload_lengths_1_14), .C(clock_c), .E(n24043), 
            .D(n174));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE i148_149 (.Q(payload_lengths_1_15), .C(clock_c), .E(n24041), 
            .D(n178));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    SB_DFFE counter_from_last_rise__i4 (.Q(counter_from_last_rise[4]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_7));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i5 (.Q(counter_from_last_rise_c[5]), .C(clock_c), 
            .E(VCC_net), .D(n23689));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i7734_3_lut_4_lut (.I0(n984), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1202), .O(n11844));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7734_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE counter_from_last_rise__i6 (.Q(\counter_from_last_rise[6] ), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_8));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i7 (.Q(\counter_from_last_rise[7] ), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_9));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i8 (.Q(\counter_from_last_rise[8] ), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_10));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i9 (.Q(\counter_from_last_rise[9] ), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_11));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i10 (.Q(\counter_from_last_rise[10] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_12));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i11 (.Q(\counter_from_last_rise[11] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_13));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i12 (.Q(\counter_from_last_rise[12] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_14));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i13 (.Q(counter_from_last_rise[13]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_15));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i14 (.Q(counter_from_last_rise[14]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_16));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i15 (.Q(counter_from_last_rise[15]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_17));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i16 (.Q(counter_from_last_rise[16]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_18));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i17 (.Q(counter_from_last_rise[17]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_19));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i18 (.Q(counter_from_last_rise[18]), .C(clock_c), 
            .E(VCC_net), .D(n8_adj_20));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i19 (.Q(\counter_from_last_rise[19] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_21));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i20 (.Q(\counter_from_last_rise[20] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_22));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i21 (.Q(\counter_from_last_rise[21] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_23));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i22 (.Q(\counter_from_last_rise[22] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_24));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i23 (.Q(\counter_from_last_rise[23] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_25));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i24 (.Q(\counter_from_last_rise[24] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_26));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i25 (.Q(\counter_from_last_rise[25] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_27));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i26 (.Q(\counter_from_last_rise[26] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_28));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i27 (.Q(\counter_from_last_rise[27] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_29));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i28 (.Q(\counter_from_last_rise[28] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_30));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i29 (.Q(\counter_from_last_rise[29] ), 
            .C(clock_c), .E(VCC_net), .D(n8_adj_31));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i30 (.Q(\counter_from_last_rise[30] ), 
            .C(clock_c), .E(VCC_net), .D(n23407));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFE counter_from_last_rise__i31 (.Q(\counter_from_last_rise[31] ), 
            .C(clock_c), .E(VCC_net), .D(n23397));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF i663__i264 (.Q(\ootx_payload_o[0][263] ), .C(clock_c), .D(n12201));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i263 (.Q(\ootx_payload_o[0][262] ), .C(clock_c), .D(n12200));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i262 (.Q(\ootx_payload_o[0][261] ), .C(clock_c), .D(n12199));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i261 (.Q(\ootx_payload_o[0][260] ), .C(clock_c), .D(n12198));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i260 (.Q(\ootx_payload_o[0][259] ), .C(clock_c), .D(n12197));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i259 (.Q(\ootx_payload_o[0][258] ), .C(clock_c), .D(n12196));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i258 (.Q(\ootx_payload_o[0][257] ), .C(clock_c), .D(n12195));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i257 (.Q(\ootx_payload_o[0][256] ), .C(clock_c), .D(n12194));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i256 (.Q(\ootx_payload_o[0][255] ), .C(clock_c), .D(n12193));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i255 (.Q(\ootx_payload_o[0][254] ), .C(clock_c), .D(n12192));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i254 (.Q(\ootx_payload_o[0][253] ), .C(clock_c), .D(n12191));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i253 (.Q(\ootx_payload_o[0][252] ), .C(clock_c), .D(n12190));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i252 (.Q(\ootx_payload_o[0][251] ), .C(clock_c), .D(n12189));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i251 (.Q(\ootx_payload_o[0][250] ), .C(clock_c), .D(n12188));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i250 (.Q(\ootx_payload_o[0][249] ), .C(clock_c), .D(n12187));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i249 (.Q(\ootx_payload_o[0][248] ), .C(clock_c), .D(n12186));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i248 (.Q(\ootx_payload_o[0][247] ), .C(clock_c), .D(n12185));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i247 (.Q(\ootx_payload_o[0][246] ), .C(clock_c), .D(n12184));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i246 (.Q(\ootx_payload_o[0][245] ), .C(clock_c), .D(n12183));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i245 (.Q(\ootx_payload_o[0][244] ), .C(clock_c), .D(n12182));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i244 (.Q(\ootx_payload_o[0][243] ), .C(clock_c), .D(n12181));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i243 (.Q(\ootx_payload_o[0][242] ), .C(clock_c), .D(n12180));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i242 (.Q(\ootx_payload_o[0][241] ), .C(clock_c), .D(n12179));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i241 (.Q(\ootx_payload_o[0][240] ), .C(clock_c), .D(n12178));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i240 (.Q(\ootx_payload_o[0][239] ), .C(clock_c), .D(n12177));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i239 (.Q(\ootx_payload_o[0][238] ), .C(clock_c), .D(n12176));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i238 (.Q(\ootx_payload_o[0][237] ), .C(clock_c), .D(n12175));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i237 (.Q(\ootx_payload_o[0][236] ), .C(clock_c), .D(n12174));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i236 (.Q(\ootx_payload_o[0][235] ), .C(clock_c), .D(n12173));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i235 (.Q(\ootx_payload_o[0][234] ), .C(clock_c), .D(n12172));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i234 (.Q(\ootx_payload_o[0][233] ), .C(clock_c), .D(n12171));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i233 (.Q(\ootx_payload_o[0][232] ), .C(clock_c), .D(n12170));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i232 (.Q(\ootx_payload_o[0][231] ), .C(clock_c), .D(n12169));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i231 (.Q(\ootx_payload_o[0][230] ), .C(clock_c), .D(n12168));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i230 (.Q(\ootx_payload_o[0][229] ), .C(clock_c), .D(n12167));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i229 (.Q(\ootx_payload_o[0][228] ), .C(clock_c), .D(n12166));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i228 (.Q(\ootx_payload_o[0][227] ), .C(clock_c), .D(n12165));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i227 (.Q(\ootx_payload_o[0][226] ), .C(clock_c), .D(n12164));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i226 (.Q(\ootx_payload_o[0][225] ), .C(clock_c), .D(n12163));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i225 (.Q(\ootx_payload_o[0][224] ), .C(clock_c), .D(n12162));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i224 (.Q(\ootx_payload_o[0][223] ), .C(clock_c), .D(n12161));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i223 (.Q(\ootx_payload_o[0][222] ), .C(clock_c), .D(n12160));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i222 (.Q(\ootx_payload_o[0][221] ), .C(clock_c), .D(n12159));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i221 (.Q(\ootx_payload_o[0][220] ), .C(clock_c), .D(n12158));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i220 (.Q(\ootx_payload_o[0][219] ), .C(clock_c), .D(n12157));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i219 (.Q(\ootx_payload_o[0][218] ), .C(clock_c), .D(n12156));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i218 (.Q(\ootx_payload_o[0][217] ), .C(clock_c), .D(n12155));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i217 (.Q(\ootx_payload_o[0][216] ), .C(clock_c), .D(n12154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i216 (.Q(\ootx_payload_o[0][215] ), .C(clock_c), .D(n12153));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i215 (.Q(\ootx_payload_o[0][214] ), .C(clock_c), .D(n12152));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i214 (.Q(\ootx_payload_o[0][213] ), .C(clock_c), .D(n12151));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i213 (.Q(\ootx_payload_o[0][212] ), .C(clock_c), .D(n12150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i212 (.Q(\ootx_payload_o[0][211] ), .C(clock_c), .D(n12149));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i211 (.Q(\ootx_payload_o[0][210] ), .C(clock_c), .D(n12148));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i210 (.Q(\ootx_payload_o[0][209] ), .C(clock_c), .D(n12147));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i209 (.Q(\ootx_payload_o[0][208] ), .C(clock_c), .D(n12146));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i208 (.Q(\ootx_payload_o[0][207] ), .C(clock_c), .D(n12145));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i207 (.Q(\ootx_payload_o[0][206] ), .C(clock_c), .D(n12144));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i206 (.Q(\ootx_payload_o[0][205] ), .C(clock_c), .D(n12143));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i205 (.Q(\ootx_payload_o[0][204] ), .C(clock_c), .D(n12142));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i204 (.Q(\ootx_payload_o[0][203] ), .C(clock_c), .D(n12141));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i203 (.Q(\ootx_payload_o[0][202] ), .C(clock_c), .D(n12140));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i202 (.Q(\ootx_payload_o[0][201] ), .C(clock_c), .D(n12139));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i201 (.Q(\ootx_payload_o[0][200] ), .C(clock_c), .D(n12138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i200 (.Q(\ootx_payload_o[0][199] ), .C(clock_c), .D(n12137));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i199 (.Q(\ootx_payload_o[0][198] ), .C(clock_c), .D(n12136));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i198 (.Q(\ootx_payload_o[0][197] ), .C(clock_c), .D(n12135));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i197 (.Q(\ootx_payload_o[0][196] ), .C(clock_c), .D(n12134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i196 (.Q(\ootx_payload_o[0][195] ), .C(clock_c), .D(n12133));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i195 (.Q(\ootx_payload_o[0][194] ), .C(clock_c), .D(n12132));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i194 (.Q(\ootx_payload_o[0][193] ), .C(clock_c), .D(n12131));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i193 (.Q(\ootx_payload_o[0][192] ), .C(clock_c), .D(n12130));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i192 (.Q(\ootx_payload_o[0][191] ), .C(clock_c), .D(n12129));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i191 (.Q(\ootx_payload_o[0][190] ), .C(clock_c), .D(n12128));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i190 (.Q(\ootx_payload_o[0][189] ), .C(clock_c), .D(n12127));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i189 (.Q(\ootx_payload_o[0][188] ), .C(clock_c), .D(n12126));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i188 (.Q(\ootx_payload_o[0][187] ), .C(clock_c), .D(n12125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i187 (.Q(\ootx_payload_o[0][186] ), .C(clock_c), .D(n12124));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i186 (.Q(\ootx_payload_o[0][185] ), .C(clock_c), .D(n12123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i185 (.Q(\ootx_payload_o[0][184] ), .C(clock_c), .D(n12122));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i184 (.Q(\ootx_payload_o[0][183] ), .C(clock_c), .D(n12121));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i183 (.Q(\ootx_payload_o[0][182] ), .C(clock_c), .D(n12120));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i182 (.Q(\ootx_payload_o[0][181] ), .C(clock_c), .D(n12119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i181 (.Q(\ootx_payload_o[0][180] ), .C(clock_c), .D(n12118));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i180 (.Q(\ootx_payload_o[0][179] ), .C(clock_c), .D(n12117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i179 (.Q(\ootx_payload_o[0][178] ), .C(clock_c), .D(n12116));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i178 (.Q(\ootx_payload_o[0][177] ), .C(clock_c), .D(n12115));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i177 (.Q(\ootx_payload_o[0][176] ), .C(clock_c), .D(n12114));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i176 (.Q(\ootx_payload_o[0][175] ), .C(clock_c), .D(n12113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i175 (.Q(\ootx_payload_o[0][174] ), .C(clock_c), .D(n12112));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i174 (.Q(\ootx_payload_o[0][173] ), .C(clock_c), .D(n12111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i173 (.Q(\ootx_payload_o[0][172] ), .C(clock_c), .D(n12110));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i172 (.Q(\ootx_payload_o[0][171] ), .C(clock_c), .D(n12109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i171 (.Q(\ootx_payload_o[0][170] ), .C(clock_c), .D(n12108));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i170 (.Q(\ootx_payload_o[0][169] ), .C(clock_c), .D(n12107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i169 (.Q(\ootx_payload_o[0][168] ), .C(clock_c), .D(n12106));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i168 (.Q(\ootx_payload_o[0][167] ), .C(clock_c), .D(n12105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i167 (.Q(\ootx_payload_o[0][166] ), .C(clock_c), .D(n12104));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i166 (.Q(\ootx_payload_o[0][165] ), .C(clock_c), .D(n12103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i165 (.Q(\ootx_payload_o[0][164] ), .C(clock_c), .D(n12102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i164 (.Q(\ootx_payload_o[0][163] ), .C(clock_c), .D(n12101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i163 (.Q(\ootx_payload_o[0][162] ), .C(clock_c), .D(n12100));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i162 (.Q(\ootx_payload_o[0][161] ), .C(clock_c), .D(n12099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i161 (.Q(\ootx_payload_o[0][160] ), .C(clock_c), .D(n12098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i160 (.Q(\ootx_payload_o[0][159] ), .C(clock_c), .D(n12097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i159 (.Q(\ootx_payload_o[0][158] ), .C(clock_c), .D(n12096));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i158 (.Q(\ootx_payload_o[0][157] ), .C(clock_c), .D(n12095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i157 (.Q(\ootx_payload_o[0][156] ), .C(clock_c), .D(n12094));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i156 (.Q(\ootx_payload_o[0][155] ), .C(clock_c), .D(n12093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i155 (.Q(\ootx_payload_o[0][154] ), .C(clock_c), .D(n12092));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i154 (.Q(\ootx_payload_o[0][153] ), .C(clock_c), .D(n12091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i153 (.Q(\ootx_payload_o[0][152] ), .C(clock_c), .D(n12090));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i152 (.Q(\ootx_payload_o[0][151] ), .C(clock_c), .D(n12089));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i151 (.Q(\ootx_payload_o[0][150] ), .C(clock_c), .D(n12088));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i150 (.Q(\ootx_payload_o[0][149] ), .C(clock_c), .D(n12087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i149 (.Q(\ootx_payload_o[0][148] ), .C(clock_c), .D(n12086));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i148 (.Q(\ootx_payload_o[0][147] ), .C(clock_c), .D(n12085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i147 (.Q(\ootx_payload_o[0][146] ), .C(clock_c), .D(n12084));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i146 (.Q(\ootx_payload_o[0][145] ), .C(clock_c), .D(n12083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i145 (.Q(\ootx_payload_o[0][144] ), .C(clock_c), .D(n12082));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i144 (.Q(\ootx_payload_o[0][143] ), .C(clock_c), .D(n12081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i143 (.Q(\ootx_payload_o[0][142] ), .C(clock_c), .D(n12080));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i142 (.Q(\ootx_payload_o[0][141] ), .C(clock_c), .D(n12079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i141 (.Q(\ootx_payload_o[0][140] ), .C(clock_c), .D(n12078));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i140 (.Q(\ootx_payload_o[0][139] ), .C(clock_c), .D(n12077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i139 (.Q(\ootx_payload_o[0][138] ), .C(clock_c), .D(n12076));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i138 (.Q(\ootx_payload_o[0][137] ), .C(clock_c), .D(n12075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i137 (.Q(\ootx_payload_o[0][136] ), .C(clock_c), .D(n12074));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i136 (.Q(\ootx_payload_o[0][135] ), .C(clock_c), .D(n12073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i135 (.Q(\ootx_payload_o[0][134] ), .C(clock_c), .D(n12072));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i134 (.Q(\ootx_payload_o[0][133] ), .C(clock_c), .D(n12071));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i133 (.Q(\ootx_payload_o[0][132] ), .C(clock_c), .D(n12070));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i132 (.Q(\ootx_payload_o[0][131] ), .C(clock_c), .D(n12069));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i131 (.Q(\ootx_payload_o[0][130] ), .C(clock_c), .D(n12068));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i130 (.Q(\ootx_payload_o[0][129] ), .C(clock_c), .D(n12067));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i129 (.Q(\ootx_payload_o[0][128] ), .C(clock_c), .D(n12066));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i128 (.Q(\ootx_payload_o[0][127] ), .C(clock_c), .D(n12065));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i127 (.Q(\ootx_payload_o[0][126] ), .C(clock_c), .D(n12064));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i126 (.Q(\ootx_payload_o[0][125] ), .C(clock_c), .D(n12063));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i125 (.Q(\ootx_payload_o[0][124] ), .C(clock_c), .D(n12062));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i124 (.Q(\ootx_payload_o[0][123] ), .C(clock_c), .D(n12061));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i123 (.Q(\ootx_payload_o[0][122] ), .C(clock_c), .D(n12060));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i122 (.Q(\ootx_payload_o[0][121] ), .C(clock_c), .D(n12059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i121 (.Q(\ootx_payload_o[0][120] ), .C(clock_c), .D(n12058));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i120 (.Q(\ootx_payload_o[0][119] ), .C(clock_c), .D(n12057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i119 (.Q(\ootx_payload_o[0][118] ), .C(clock_c), .D(n12056));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i118 (.Q(\ootx_payload_o[0][117] ), .C(clock_c), .D(n12055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i117 (.Q(\ootx_payload_o[0][116] ), .C(clock_c), .D(n12054));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i116 (.Q(\ootx_payload_o[0][115] ), .C(clock_c), .D(n12053));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i115 (.Q(\ootx_payload_o[0][114] ), .C(clock_c), .D(n12052));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i114 (.Q(\ootx_payload_o[0][113] ), .C(clock_c), .D(n12051));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i113 (.Q(\ootx_payload_o[0][112] ), .C(clock_c), .D(n12050));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i112 (.Q(\ootx_payload_o[0][111] ), .C(clock_c), .D(n12049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i111 (.Q(\ootx_payload_o[0][110] ), .C(clock_c), .D(n12048));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i110 (.Q(\ootx_payload_o[0][109] ), .C(clock_c), .D(n12047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i109 (.Q(\ootx_payload_o[0][108] ), .C(clock_c), .D(n12046));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i108 (.Q(\ootx_payload_o[0][107] ), .C(clock_c), .D(n12045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i107 (.Q(\ootx_payload_o[0][106] ), .C(clock_c), .D(n12044));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i106 (.Q(\ootx_payload_o[0][105] ), .C(clock_c), .D(n12043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i105 (.Q(\ootx_payload_o[0][104] ), .C(clock_c), .D(n12042));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i104 (.Q(\ootx_payload_o[0][103] ), .C(clock_c), .D(n12041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i103 (.Q(\ootx_payload_o[0][102] ), .C(clock_c), .D(n12040));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i102 (.Q(\ootx_payload_o[0][101] ), .C(clock_c), .D(n12039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i101 (.Q(\ootx_payload_o[0][100] ), .C(clock_c), .D(n12038));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i100 (.Q(\ootx_payload_o[0][99] ), .C(clock_c), .D(n12037));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i99 (.Q(\ootx_payload_o[0][98] ), .C(clock_c), .D(n12036));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i98 (.Q(\ootx_payload_o[0][97] ), .C(clock_c), .D(n12035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i97 (.Q(\ootx_payload_o[0][96] ), .C(clock_c), .D(n12034));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i96 (.Q(\ootx_payload_o[0][95] ), .C(clock_c), .D(n12033));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i95 (.Q(\ootx_payload_o[0][94] ), .C(clock_c), .D(n12032));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i94 (.Q(\ootx_payload_o[0][93] ), .C(clock_c), .D(n12031));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i93 (.Q(\ootx_payload_o[0][92] ), .C(clock_c), .D(n12030));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i92 (.Q(\ootx_payload_o[0][91] ), .C(clock_c), .D(n12029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i91 (.Q(\ootx_payload_o[0][90] ), .C(clock_c), .D(n12028));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i90 (.Q(\ootx_payload_o[0][89] ), .C(clock_c), .D(n12027));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i89 (.Q(\ootx_payload_o[0][88] ), .C(clock_c), .D(n12026));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i88 (.Q(\ootx_payload_o[0][87] ), .C(clock_c), .D(n12025));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i87 (.Q(\ootx_payload_o[0][86] ), .C(clock_c), .D(n12024));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i86 (.Q(\ootx_payload_o[0][85] ), .C(clock_c), .D(n12023));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i85 (.Q(\ootx_payload_o[0][84] ), .C(clock_c), .D(n12022));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i84 (.Q(\ootx_payload_o[0][83] ), .C(clock_c), .D(n12021));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i83 (.Q(\ootx_payload_o[0][82] ), .C(clock_c), .D(n12020));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i82 (.Q(\ootx_payload_o[0][81] ), .C(clock_c), .D(n12019));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i81 (.Q(\ootx_payload_o[0][80] ), .C(clock_c), .D(n12018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i80 (.Q(\ootx_payload_o[0][79] ), .C(clock_c), .D(n12017));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i79 (.Q(\ootx_payload_o[0][78] ), .C(clock_c), .D(n12016));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i78 (.Q(\ootx_payload_o[0][77] ), .C(clock_c), .D(n12015));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i77 (.Q(\ootx_payload_o[0][76] ), .C(clock_c), .D(n12014));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i76 (.Q(\ootx_payload_o[0][75] ), .C(clock_c), .D(n12013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i75 (.Q(\ootx_payload_o[0][74] ), .C(clock_c), .D(n12012));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i74 (.Q(\ootx_payload_o[0][73] ), .C(clock_c), .D(n12011));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i73 (.Q(\ootx_payload_o[0][72] ), .C(clock_c), .D(n12010));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i72 (.Q(\ootx_payload_o[0][71] ), .C(clock_c), .D(n12009));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i71 (.Q(\ootx_payload_o[0][70] ), .C(clock_c), .D(n12008));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i70 (.Q(\ootx_payload_o[0][69] ), .C(clock_c), .D(n12007));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i69 (.Q(\ootx_payload_o[0][68] ), .C(clock_c), .D(n12006));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i68 (.Q(\ootx_payload_o[0][67] ), .C(clock_c), .D(n12005));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i67 (.Q(\ootx_payload_o[0][66] ), .C(clock_c), .D(n12004));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i66 (.Q(\ootx_payload_o[0][65] ), .C(clock_c), .D(n12003));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i65 (.Q(\ootx_payload_o[0][64] ), .C(clock_c), .D(n12002));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i64 (.Q(\ootx_payload_o[0][63] ), .C(clock_c), .D(n12001));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i63 (.Q(\ootx_payload_o[0][62] ), .C(clock_c), .D(n12000));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i62 (.Q(\ootx_payload_o[0][61] ), .C(clock_c), .D(n11999));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i61 (.Q(\ootx_payload_o[0][60] ), .C(clock_c), .D(n11998));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i60 (.Q(\ootx_payload_o[0][59] ), .C(clock_c), .D(n11997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i59 (.Q(\ootx_payload_o[0][58] ), .C(clock_c), .D(n11996));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i58 (.Q(\ootx_payload_o[0][57] ), .C(clock_c), .D(n11995));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i57 (.Q(\ootx_payload_o[0][56] ), .C(clock_c), .D(n11994));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i56 (.Q(\ootx_payload_o[0][55] ), .C(clock_c), .D(n11993));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i55 (.Q(\ootx_payload_o[0][54] ), .C(clock_c), .D(n11992));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i54 (.Q(\ootx_payload_o[0][53] ), .C(clock_c), .D(n11991));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i53 (.Q(\ootx_payload_o[0][52] ), .C(clock_c), .D(n11990));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFFER ootx_states_1__i0_i1 (.Q(\ootx_states[1] [1]), .C(clock_c), 
            .E(n23147), .D(ootx_states_1__1__N_896[1]), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF i560_561 (.Q(ootx_payloads_0_94), .C(clock_c), .D(n11115));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_4_lut (.I0(\lighthouse[0] ), .I1(ootx_payloads_N_1744[0]), 
            .I2(n31), .I3(n22_adj_1846), .O(n34_c));
    defparam i1_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 i7142_3_lut_4_lut (.I0(n984), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_231), .O(n11252));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7142_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7711_3_lut_4_lut (.I0(n938), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1225), .O(n11821));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7711_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_49 (.I0(n83), .I1(n19313), .I2(n2851[30]), .I3(n60_c), 
            .O(n608_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i1_4_lut_adj_49.LUT_INIT = 16'h222a;
    SB_DFF i663__i52 (.Q(\ootx_payload_o[0][51] ), .C(clock_c), .D(n11989));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 i3_4_lut_adj_50 (.I0(n2851[27]), .I1(n2851[28]), .I2(n2851[29]), 
            .I3(n2851[30]), .O(n19313));
    defparam i3_4_lut_adj_50.LUT_INIT = 16'hfffe;
    SB_DFF i663__i51 (.Q(\ootx_payload_o[0][50] ), .C(clock_c), .D(n11988));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 i1_4_lut_adj_51 (.I0(new_data), .I1(ootx_payloads_N_1744[1]), 
            .I2(n34_c), .I3(n27), .O(n23163));
    defparam i1_4_lut_adj_51.LUT_INIT = 16'ha2a0;
    SB_LUT4 mod_155_add_2009_25_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n22777), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i663__i50 (.Q(\ootx_payload_o[0][49] ), .C(clock_c), .D(n11987));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_CARRY add_154_16 (.CI(n22257), .I0(n2849[14]), .I1(GND_net), .CO(n22258));
    SB_DFF i663__i49 (.Q(\ootx_payload_o[0][48] ), .C(clock_c), .D(n11986));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i48 (.Q(\ootx_payload_o[0][47] ), .C(clock_c), .D(n11985));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_CARRY mod_155_add_1942_19 (.CI(n22744), .I0(n2796), .I1(n2819), 
            .CO(n22745));
    SB_LUT4 add_355_14_lut (.I0(GND_net), .I1(\counter_from_last_rise[12] ), 
            .I2(GND_net), .I3(n22286), .O(n6333[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF i663__i47 (.Q(\ootx_payload_o[0][46] ), .C(clock_c), .D(n11984));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i46 (.Q(\ootx_payload_o[0][45] ), .C(clock_c), .D(n11983));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 add_154_15_lut (.I0(GND_net), .I1(n2849[13]), .I2(GND_net), 
            .I3(n22256), .O(n2851[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7721_3_lut_4_lut (.I0(n958), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1215), .O(n11831));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7721_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i663__i45 (.Q(\ootx_payload_o[0][44] ), .C(clock_c), .D(n11982));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_CARRY mod_155_add_2076_29 (.CI(n22809), .I0(n2986), .I1(n3017), 
            .CO(n22810));
    SB_LUT4 mod_155_add_1808_15_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n22689), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_18_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[16]), 
            .I2(GND_net), .I3(n22229), .O(n337[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1330_2_lut (.I0(n2851[28]), .I1(n2851[27]), .I2(GND_net), 
            .I3(GND_net), .O(n58_adj_1820));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i1330_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_155_add_1540_7 (.CI(n22591), .I0(n2208), .I1(n2225), 
            .CO(n22592));
    SB_CARRY add_66_18 (.CI(n22229), .I0(ootx_payloads_N_1699[16]), .I1(GND_net), 
            .CO(n22230));
    SB_LUT4 mux_431_Mux_1_i3_4_lut (.I0(n10802), .I1(n30), .I2(ootx_payloads_N_1744[1]), 
            .I3(\lighthouse[0] ), .O(ootx_states_0__1__N_898[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[6] 189[13])
    defparam mux_431_Mux_1_i3_4_lut.LUT_INIT = 16'h303a;
    SB_CARRY mod_155_add_2009_25 (.CI(n22777), .I0(n2890), .I1(n2918), 
            .CO(n22778));
    SB_DFF i663__i44 (.Q(\ootx_payload_o[0][43] ), .C(clock_c), .D(n11981));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 i7129_3_lut_4_lut (.I0(n958), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_218), .O(n11239));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7129_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1004_15_lut (.I0(n1400_c), .I1(n1400_c), .I2(n1433_c), 
            .I3(n22467), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_15 (.CI(n22256), .I0(n2849[13]), .I1(GND_net), .CO(n22257));
    SB_DFF i663__i43 (.Q(\ootx_payload_o[0][42] ), .C(clock_c), .D(n11980));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 mod_155_add_1540_6_lut (.I0(n2209), .I1(n2209), .I2(n25179), 
            .I3(n22590), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1004_14_lut (.I0(n1401_c), .I1(n1401_c), .I2(n1433_c), 
            .I3(n22466), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_14_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i663__i42 (.Q(\ootx_payload_o[0][41] ), .C(clock_c), .D(n11979));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i41 (.Q(\ootx_payload_o[0][40] ), .C(clock_c), .D(n11978));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_CARRY mod_155_add_1808_15 (.CI(n22689), .I0(n2600), .I1(n2621), 
            .CO(n22690));
    SB_DFF i663__i40 (.Q(\ootx_payload_o[0][39] ), .C(clock_c), .D(n11977));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 mod_155_add_1808_14_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n22688), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1540_6 (.CI(n22590), .I0(n2209), .I1(n25179), 
            .CO(n22591));
    SB_LUT4 i7733_3_lut_4_lut (.I0(n982), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1203), .O(n11843));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7733_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1004_14 (.CI(n22466), .I0(n1401_c), .I1(n1433_c), 
            .CO(n22467));
    SB_LUT4 i7141_3_lut_4_lut (.I0(n982), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_230), .O(n11251));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7141_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i663__i39 (.Q(\ootx_payload_o[0][38] ), .C(clock_c), .D(n11976));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i557_558 (.Q(ootx_payloads_0_93), .C(clock_c), .D(n11114));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i663__i38 (.Q(\ootx_payload_o[0][37] ), .C(clock_c), .D(n11975));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 i7119_3_lut_4_lut (.I0(n938), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_208), .O(n11229));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7119_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_52 (.I0(n2851[26]), .I1(n612_c), .I2(n611), .I3(n610_c), 
            .O(n22887));
    defparam i3_4_lut_adj_52.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1540_5_lut (.I0(n2210), .I1(n2210), .I2(n2225), 
            .I3(n22589), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i663__i37 (.Q(\ootx_payload_o[0][36] ), .C(clock_c), .D(n11974));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 mod_155_add_1004_13_lut (.I0(n1402_c), .I1(n1402_c), .I2(n1433_c), 
            .I3(n22465), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_14 (.CI(n22286), .I0(\counter_from_last_rise[12] ), 
            .I1(GND_net), .CO(n22287));
    SB_LUT4 i15377_3_lut (.I0(n22887), .I1(n608_c), .I2(n609), .I3(GND_net), 
            .O(n641));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i15377_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_155_i474_3_lut (.I0(n612_c), .I1(n89[27]), .I2(n641), 
            .I3(GND_net), .O(n711));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_i475_3_lut (.I0(n2851[26]), .I1(n89[26]), .I2(n641), 
            .I3(GND_net), .O(n712_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1942_18_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n22743), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_14_lut (.I0(GND_net), .I1(n2849[12]), .I2(GND_net), 
            .I3(n22255), .O(n2851[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1808_14 (.CI(n22688), .I0(n2601), .I1(n2621), 
            .CO(n22689));
    SB_CARRY add_154_14 (.CI(n22255), .I0(n2849[12]), .I1(GND_net), .CO(n22256));
    SB_LUT4 mod_155_add_1808_13_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n22687), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i663__i36 (.Q(\ootx_payload_o[0][35] ), .C(clock_c), .D(n11973));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF sensor_state_482 (.Q(sensor_state), .C(clock_c), .D(n23693));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF i663__i35 (.Q(\ootx_payload_o[0][34] ), .C(clock_c), .D(n11972));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i34 (.Q(\ootx_payload_o[0][33] ), .C(clock_c), .D(n11971));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i33 (.Q(\ootx_payload_o[0][32] ), .C(clock_c), .D(n11970));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 add_355_13_lut (.I0(GND_net), .I1(\counter_from_last_rise[11] ), 
            .I2(GND_net), .I3(n22285), .O(n6333[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF i663__i32 (.Q(\ootx_payload_o[0][31] ), .C(clock_c), .D(n11969));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i31 (.Q(\ootx_payload_o[0][30] ), .C(clock_c), .D(n11968));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 i3_4_lut_adj_53 (.I0(n2851[25]), .I1(n712_c), .I2(n711), .I3(n710_c), 
            .O(n22886));
    defparam i3_4_lut_adj_53.LUT_INIT = 16'hfffe;
    SB_DFF i663__i30 (.Q(\ootx_payload_o[0][29] ), .C(clock_c), .D(n11967));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i29 (.Q(\ootx_payload_o[0][28] ), .C(clock_c), .D(n11966));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i28 (.Q(\ootx_payload_o[0][27] ), .C(clock_c), .D(n11965));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i27 (.Q(\ootx_payload_o[0][26] ), .C(clock_c), .D(n11964));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 i19432_4_lut (.I0(n707), .I1(n22886), .I2(n708_c), .I3(n709), 
            .O(n740_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i19432_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 add_154_13_lut (.I0(GND_net), .I1(n2849[11]), .I2(GND_net), 
            .I3(n22254), .O(n2851[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF i663__i26 (.Q(\ootx_payload_o[0][25] ), .C(clock_c), .D(n11963));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i25 (.Q(\ootx_payload_o[0][24] ), .C(clock_c), .D(n11962));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_CARRY mod_155_add_1540_5 (.CI(n22589), .I0(n2210), .I1(n2225), 
            .CO(n22590));
    SB_DFF i663__i24 (.Q(\ootx_payload_o[0][23] ), .C(clock_c), .D(n11961));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i23 (.Q(\ootx_payload_o[0][22] ), .C(clock_c), .D(n11960));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 mod_155_i473_3_lut (.I0(n611), .I1(n89[28]), .I2(n641), .I3(GND_net), 
            .O(n710_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i473_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i663__i22 (.Q(\ootx_payload_o[0][21] ), .C(clock_c), .D(n11959));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i554_555 (.Q(ootx_payloads_0_92), .C(clock_c), .D(n11113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i6990_3_lut_4_lut (.I0(n680), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_79), .O(n11100));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6990_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_i540_3_lut (.I0(n710_c), .I1(n773[28]), .I2(n740_c), 
            .I3(GND_net), .O(n809));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam mod_155_i540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7582_3_lut_4_lut (.I0(n680), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1354), .O(n11692));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7582_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_54 (.I0(n806_c), .I1(n807), .I2(n808_c), .I3(GND_net), 
            .O(n23950));
    defparam i2_3_lut_adj_54.LUT_INIT = 16'hfefe;
    SB_LUT4 i7006_3_lut_4_lut (.I0(n712), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_95), .O(n11116));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7006_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut (.I0(n812_c), .I1(n810_c), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_55 (.I0(n29_adj_1850), .I1(n23950), .I2(n809), 
            .I3(n6), .O(n839));
    defparam i1_4_lut_adj_55.LUT_INIT = 16'hfcec;
    SB_LUT4 i7598_3_lut_4_lut (.I0(n712), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1338), .O(n11708));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7598_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut (.I0(n2851[24]), .I1(n811), .I2(GND_net), .I3(GND_net), 
            .O(n29_adj_1850));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20353_2_lut (.I0(n71[26]), .I1(n71[24]), .I2(GND_net), .I3(GND_net), 
            .O(n24713));
    defparam i20353_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20460_4_lut (.I0(n71[30]), .I1(n71[28]), .I2(n71[31]), .I3(n71[29]), 
            .O(n24553));
    defparam i20460_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_56 (.I0(n29_adj_1850), .I1(n2851[23]), .I2(n24713), 
            .I3(n839), .O(n4_adj_1851));
    defparam i1_4_lut_adj_56.LUT_INIT = 16'hfcee;
    SB_LUT4 i34_4_lut (.I0(n23950), .I1(n24553), .I2(n839), .I3(n809), 
            .O(n39_c));
    defparam i34_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i15280_4_lut (.I0(n911), .I1(n39_c), .I2(n909), .I3(n4_adj_1851), 
            .O(n938_c));
    defparam i15280_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i9431_3_lut (.I0(n806_c), .I1(n71[31]), .I2(n839), .I3(GND_net), 
            .O(n905));
    defparam i9431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i126_2_lut_3_lut (.I0(n29_adj_1852), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n126_adj_1853));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i126_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i125_2_lut_3_lut (.I0(n29_adj_1852), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i125_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i30_2_lut_3_lut (.I0(n13_adj_1854), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(GND_net), .O(n30_adj_1855));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i30_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i29_2_lut_3_lut (.I0(n13_adj_1854), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(GND_net), .O(n29_adj_1852));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i29_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 Mux_16_i1_3_lut (.I0(bit_counters_0_20), .I1(bit_counters_1_20), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[20]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_16_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20525_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25193));
    defparam i20525_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_57 (.I0(n2851[8]), .I1(n2412), .I2(n2411), .I3(n2410), 
            .O(n22896));
    defparam i3_4_lut_adj_57.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n2408), .I1(n22896), .I2(n2409), .I3(GND_net), 
            .O(n23));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i11_4_lut_adj_58 (.I0(n2404), .I1(n2403), .I2(n2407), .I3(n2398), 
            .O(n31_adj_1856));
    defparam i11_4_lut_adj_58.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(counter_from_last_rise_c[5]), .I1(n24697), .I2(n2282), 
            .I3(n6333_c[5]), .O(n23689));
    defparam i18_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i16_4_lut_adj_59 (.I0(n31_adj_1856), .I1(n23), .I2(n2399), 
            .I3(n2392), .O(n36));
    defparam i16_4_lut_adj_59.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2391), .I1(n2394), .I2(n2393), .I3(n2402), 
            .O(n34_adj_1857));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_60 (.I0(n2390), .I1(n2400), .I2(n2396), .I3(n2405), 
            .O(n35_adj_1858));
    defparam i15_4_lut_adj_60.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_61 (.I0(n2406), .I1(n2397), .I2(n2395), .I3(n2401), 
            .O(n33));
    defparam i13_4_lut_adj_61.LUT_INIT = 16'hfffe;
    SB_LUT4 add_66_17_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[15] ), 
            .I2(GND_net), .I3(n22228), .O(n337[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2076_28_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n22808), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1004_13 (.CI(n22465), .I0(n1402_c), .I1(n1433_c), 
            .CO(n22466));
    SB_LUT4 i19_4_lut (.I0(n33), .I1(n35_adj_1858), .I2(n34_adj_1857), 
            .I3(n36), .O(n2423));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 Mux_15_i1_3_lut (.I0(bit_counters_0_21), .I1(bit_counters_1_21), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[21]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(n1005), .I1(n1006_c), .I2(n1008_c), .I3(n1004_c), 
            .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 PrioSelect_141_i2_3_lut (.I0(data), .I1(n4485[14]), .I2(n34[1]), 
            .I3(GND_net), .O(n174));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_141_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_62 (.I0(n2851[22]), .I1(n1012_c), .I2(n1011), 
            .I3(n1010_c), .O(n22876));
    defparam i3_4_lut_adj_62.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(n22876), .I1(n10), .I2(n1007), .I3(n1009), 
            .O(n1037));
    defparam i5_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_1_lut (.I0(reset_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2282));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i551_552 (.Q(ootx_payloads_0_91), .C(clock_c), .D(n11112));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i548_549 (.Q(ootx_payloads_0_90), .C(clock_c), .D(n11111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i545_546 (.Q(ootx_payloads_0_89), .C(clock_c), .D(n11110));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i542_543 (.Q(ootx_payloads_0_88), .C(clock_c), .D(n11109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i539_540 (.Q(ootx_payloads_0_87), .C(clock_c), .D(n11108));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i536_537 (.Q(ootx_payloads_0_86), .C(clock_c), .D(n11107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut (.I0(n38_c), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n86_adj_1860));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i86_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut (.I0(n38_c), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n85));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i85_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i533_534 (.Q(ootx_payloads_0_85), .C(clock_c), .D(n11106));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1540_4_lut (.I0(n2211), .I1(n2211), .I2(n2225), 
            .I3(n22588), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i530_531 (.Q(ootx_payloads_0_84), .C(clock_c), .D(n11105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i527_528 (.Q(ootx_payloads_0_83), .C(clock_c), .D(n11104));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 EnabledDecoder_2_i13_2_lut_3_lut (.I0(ootx_payloads_N_1685), .I1(ootx_payloads_N_1699[0]), 
            .I2(ootx_payloads_N_1699[1]), .I3(GND_net), .O(n13_adj_1854));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i13_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i524_525 (.Q(ootx_payloads_0_82), .C(clock_c), .D(n11103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i663__i21 (.Q(\ootx_payload_o[0][20] ), .C(clock_c), .D(n11958));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 mod_155_add_1004_12_lut (.I0(n1403_c), .I1(n1403_c), .I2(n1433_c), 
            .I3(n22464), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i663__i20 (.Q(\ootx_payload_o[0][19] ), .C(clock_c), .D(n11957));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 Mux_14_i1_3_lut (.I0(bit_counters_0_22), .I1(bit_counters_1_22), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[22]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_63 (.I0(n2851[13]), .I1(n1912), .I2(n1911), .I3(n1910), 
            .O(n22944));
    defparam i3_4_lut_adj_63.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_64 (.I0(n1906), .I1(n1900), .I2(n1903), .I3(n1905), 
            .O(n26_adj_1861));
    defparam i11_4_lut_adj_64.LUT_INIT = 16'hfffe;
    SB_DFF i663__i19 (.Q(\ootx_payload_o[0][18] ), .C(clock_c), .D(n11956));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i18 (.Q(\ootx_payload_o[0][17] ), .C(clock_c), .D(n11955));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i17 (.Q(\ootx_payload_o[0][16] ), .C(clock_c), .D(n11954));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i16 (.Q(\ootx_payload_o[0][15] ), .C(clock_c), .D(n11953));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i15 (.Q(\ootx_payload_o[0][14] ), .C(clock_c), .D(n11952));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i14 (.Q(\ootx_payload_o[0][13] ), .C(clock_c), .D(n11951));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i13 (.Q(\ootx_payload_o[0][12] ), .C(clock_c), .D(n11950));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i12 (.Q(\ootx_payload_o[0][11] ), .C(clock_c), .D(n11949));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i11 (.Q(\ootx_payload_o[0][10] ), .C(clock_c), .D(n11948));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i10 (.Q(\ootx_payload_o[0][9] ), .C(clock_c), .D(n11947));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i9 (.Q(\ootx_payload_o[0][8] ), .C(clock_c), .D(n11946));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i8 (.Q(\ootx_payload_o[0][7] ), .C(clock_c), .D(n11945));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i7 (.Q(\ootx_payload_o[0][6] ), .C(clock_c), .D(n11944));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i6 (.Q(\ootx_payload_o[0][5] ), .C(clock_c), .D(n11943));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i5 (.Q(\ootx_payload_o[0][4] ), .C(clock_c), .D(n11942));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i4 (.Q(\ootx_payload_o[0][3] ), .C(clock_c), .D(n11941));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i3 (.Q(\ootx_payload_o[0][2] ), .C(clock_c), .D(n11940));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF i663__i2 (.Q(\ootx_payload_o[0][1] ), .C(clock_c), .D(n11939));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_DFF ootx_crc32_2_o_i0_i31 (.Q(\ootx_crc32_o[1] [31]), .C(clock_c), 
           .D(n11938));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i30 (.Q(\ootx_crc32_o[1] [30]), .C(clock_c), 
           .D(n11937));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i29 (.Q(\ootx_crc32_o[1] [29]), .C(clock_c), 
           .D(n11936));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i28 (.Q(\ootx_crc32_o[1] [28]), .C(clock_c), 
           .D(n11935));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i27 (.Q(\ootx_crc32_o[1] [27]), .C(clock_c), 
           .D(n11934));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i26 (.Q(\ootx_crc32_o[1] [26]), .C(clock_c), 
           .D(n11933));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i25 (.Q(\ootx_crc32_o[1] [25]), .C(clock_c), 
           .D(n11932));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i24 (.Q(\ootx_crc32_o[1] [24]), .C(clock_c), 
           .D(n11931));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i23 (.Q(\ootx_crc32_o[1] [23]), .C(clock_c), 
           .D(n11930));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i22 (.Q(\ootx_crc32_o[1] [22]), .C(clock_c), 
           .D(n11929));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i21 (.Q(\ootx_crc32_o[1] [21]), .C(clock_c), 
           .D(n11928));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i20 (.Q(\ootx_crc32_o[1] [20]), .C(clock_c), 
           .D(n11927));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i19 (.Q(\ootx_crc32_o[1] [19]), .C(clock_c), 
           .D(n11926));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i9_4_lut_adj_65 (.I0(n1898), .I1(n1895), .I2(n1896), .I3(n1897), 
            .O(n24_adj_1862));
    defparam i9_4_lut_adj_65.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_66 (.I0(n1904), .I1(n1902), .I2(n1901), .I3(n1899), 
            .O(n25_c));
    defparam i10_4_lut_adj_66.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_67 (.I0(n22944), .I1(n1908), .I2(n1909), .I3(n1907), 
            .O(n23_adj_1863));
    defparam i8_4_lut_adj_67.LUT_INIT = 16'hffec;
    SB_LUT4 i14_4_lut_adj_68 (.I0(n23_adj_1863), .I1(n25_c), .I2(n24_adj_1862), 
            .I3(n26_adj_1861), .O(n1928));
    defparam i14_4_lut_adj_68.LUT_INIT = 16'hfffe;
    SB_LUT4 i20519_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25187));
    defparam i20519_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20522_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25190));
    defparam i20522_1_lut.LUT_INIT = 16'h5555;
    SB_DFF ootx_crc32_2_o_i0_i18 (.Q(\ootx_crc32_o[1] [18]), .C(clock_c), 
           .D(n11925));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i17 (.Q(\ootx_crc32_o[1] [17]), .C(clock_c), 
           .D(n11924));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i16 (.Q(\ootx_crc32_o[1] [16]), .C(clock_c), 
           .D(n11923));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i15 (.Q(\ootx_crc32_o[1] [15]), .C(clock_c), 
           .D(n11922));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i14 (.Q(\ootx_crc32_o[1] [14]), .C(clock_c), 
           .D(n11921));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i13 (.Q(\ootx_crc32_o[1] [13]), .C(clock_c), 
           .D(n11920));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i12 (.Q(\ootx_crc32_o[1] [12]), .C(clock_c), 
           .D(n11919));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i11 (.Q(\ootx_crc32_o[1] [11]), .C(clock_c), 
           .D(n11918));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i10 (.Q(\ootx_crc32_o[1] [10]), .C(clock_c), 
           .D(n11917));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i9 (.Q(\ootx_crc32_o[1] [9]), .C(clock_c), 
           .D(n11916));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i8 (.Q(\ootx_crc32_o[1] [8]), .C(clock_c), 
           .D(n11915));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i7 (.Q(\ootx_crc32_o[1] [7]), .C(clock_c), 
           .D(n11914));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i6 (.Q(\ootx_crc32_o[1] [6]), .C(clock_c), 
           .D(n11913));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i5 (.Q(\ootx_crc32_o[1] [5]), .C(clock_c), 
           .D(n11912));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i4 (.Q(\ootx_crc32_o[1] [4]), .C(clock_c), 
           .D(n11911));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i3 (.Q(\ootx_crc32_o[1] [3]), .C(clock_c), 
           .D(n11910));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i2 (.Q(\ootx_crc32_o[1] [2]), .C(clock_c), 
           .D(n11909));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_2_o_i0_i1 (.Q(\ootx_crc32_o[1] [1]), .C(clock_c), 
           .D(n11908));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i31 (.Q(\ootx_crc32_o[0] [31]), .C(clock_c), 
           .D(n11907));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i30 (.Q(\ootx_crc32_o[0] [30]), .C(clock_c), 
           .D(n11906));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i29 (.Q(\ootx_crc32_o[0] [29]), .C(clock_c), 
           .D(n11905));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i28 (.Q(\ootx_crc32_o[0] [28]), .C(clock_c), 
           .D(n11904));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i27 (.Q(\ootx_crc32_o[0] [27]), .C(clock_c), 
           .D(n11903));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i26 (.Q(\ootx_crc32_o[0] [26]), .C(clock_c), 
           .D(n11902));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i25 (.Q(\ootx_crc32_o[0] [25]), .C(clock_c), 
           .D(n11901));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i24 (.Q(\ootx_crc32_o[0] [24]), .C(clock_c), 
           .D(n11900));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i23 (.Q(\ootx_crc32_o[0] [23]), .C(clock_c), 
           .D(n11899));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 EnabledDecoder_2_i17_2_lut_3_lut_4_lut (.I0(ootx_payloads_N_1685), 
            .I1(ootx_payloads_N_1699[0]), .I2(ootx_payloads_N_1699[2]), 
            .I3(ootx_payloads_N_1699[1]), .O(n17_adj_1864));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i17_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i18_2_lut_3_lut_4_lut (.I0(ootx_payloads_N_1685), 
            .I1(ootx_payloads_N_1699[0]), .I2(ootx_payloads_N_1699[2]), 
            .I3(ootx_payloads_N_1699[1]), .O(n18_adj_1865));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i18_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_1808_13 (.CI(n22687), .I0(n2602), .I1(n2621), 
            .CO(n22688));
    SB_DFF ootx_crc32_1_o_i0_i22 (.Q(\ootx_crc32_o[0] [22]), .C(clock_c), 
           .D(n11898));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i21 (.Q(\ootx_crc32_o[0] [21]), .C(clock_c), 
           .D(n11897));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i20 (.Q(\ootx_crc32_o[0] [20]), .C(clock_c), 
           .D(n11896));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i19 (.Q(\ootx_crc32_o[0] [19]), .C(clock_c), 
           .D(n11895));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i18 (.Q(\ootx_crc32_o[0] [18]), .C(clock_c), 
           .D(n11894));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i17 (.Q(\ootx_crc32_o[0] [17]), .C(clock_c), 
           .D(n11893));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i16 (.Q(\ootx_crc32_o[0] [16]), .C(clock_c), 
           .D(n11892));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i15 (.Q(\ootx_crc32_o[0] [15]), .C(clock_c), 
           .D(n11891));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i14 (.Q(\ootx_crc32_o[0] [14]), .C(clock_c), 
           .D(n11890));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i13 (.Q(\ootx_crc32_o[0] [13]), .C(clock_c), 
           .D(n11889));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i12 (.Q(\ootx_crc32_o[0] [12]), .C(clock_c), 
           .D(n11888));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i11 (.Q(\ootx_crc32_o[0] [11]), .C(clock_c), 
           .D(n11887));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i10 (.Q(\ootx_crc32_o[0] [10]), .C(clock_c), 
           .D(n11886));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i9 (.Q(\ootx_crc32_o[0] [9]), .C(clock_c), 
           .D(n11885));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i8 (.Q(\ootx_crc32_o[0] [8]), .C(clock_c), 
           .D(n11884));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i7 (.Q(\ootx_crc32_o[0] [7]), .C(clock_c), 
           .D(n11883));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i6 (.Q(\ootx_crc32_o[0] [6]), .C(clock_c), 
           .D(n11882));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i5 (.Q(\ootx_crc32_o[0] [5]), .C(clock_c), 
           .D(n11881));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i4 (.Q(\ootx_crc32_o[0] [4]), .C(clock_c), 
           .D(n11880));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i3 (.Q(\ootx_crc32_o[0] [3]), .C(clock_c), 
           .D(n11879));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i2 (.Q(\ootx_crc32_o[0] [2]), .C(clock_c), 
           .D(n11878));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_crc32_1_o_i0_i1 (.Q(\ootx_crc32_o[0] [1]), .C(clock_c), 
           .D(n11877));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF i1067_1068 (.Q(n1170), .C(clock_c), .D(n11876));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1064_1065 (.Q(n1171), .C(clock_c), .D(n11875));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1061_1062 (.Q(n1172), .C(clock_c), .D(n11874));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1058_1059 (.Q(n1173), .C(clock_c), .D(n11873));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1055_1056 (.Q(n1174), .C(clock_c), .D(n11872));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1052_1053 (.Q(n1175), .C(clock_c), .D(n11871));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1049_1050 (.Q(n1176), .C(clock_c), .D(n11870));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1046_1047 (.Q(n1177), .C(clock_c), .D(n11869));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1043_1044 (.Q(n1178), .C(clock_c), .D(n11868));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i3_4_lut_adj_69 (.I0(n2851[5]), .I1(n2712), .I2(n2711), .I3(n2710), 
            .O(n22893));
    defparam i3_4_lut_adj_69.LUT_INIT = 16'hfffe;
    SB_DFF i1040_1041 (.Q(n1179), .C(clock_c), .D(n11867));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i13_4_lut_adj_70 (.I0(n2690), .I1(n2697), .I2(n2708), .I3(n2689), 
            .O(n36_adj_1866));
    defparam i13_4_lut_adj_70.LUT_INIT = 16'hfffe;
    SB_DFF i1037_1038 (.Q(n1180), .C(clock_c), .D(n11866));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1034_1035 (.Q(n1181), .C(clock_c), .D(n11865));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1540_4 (.CI(n22588), .I0(n2211), .I1(n2225), 
            .CO(n22589));
    SB_DFF i1031_1032 (.Q(n1182), .C(clock_c), .D(n11864));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1004_12 (.CI(n22464), .I0(n1403_c), .I1(n1433_c), 
            .CO(n22465));
    SB_DFF i1028_1029 (.Q(n1183), .C(clock_c), .D(n11863));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1025_1026 (.Q(n1184), .C(clock_c), .D(n11862));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i9_3_lut_adj_71 (.I0(n22893), .I1(n2703), .I2(n2709), .I3(GND_net), 
            .O(n32_adj_1867));
    defparam i9_3_lut_adj_71.LUT_INIT = 16'hecec;
    SB_DFF i1022_1023 (.Q(n1185), .C(clock_c), .D(n11861));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1019_1020 (.Q(n1186), .C(clock_c), .D(n11860));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i17_4_lut (.I0(n2706), .I1(n2707), .I2(n2704), .I3(n2705), 
            .O(n40_c));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF i1016_1017 (.Q(n1187), .C(clock_c), .D(n11859));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1013_1014 (.Q(n1188), .C(clock_c), .D(n11858));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i15_4_lut_adj_72 (.I0(n2701), .I1(n2696), .I2(n2695), .I3(n2688), 
            .O(n38_adj_1868));
    defparam i15_4_lut_adj_72.LUT_INIT = 16'hfffe;
    SB_DFF i1010_1011 (.Q(n1189), .C(clock_c), .D(n11857));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1007_1008 (.Q(n1190), .C(clock_c), .D(n11856));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i521_522 (.Q(ootx_payloads_0_81), .C(clock_c), .D(n11102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i14_4_lut_adj_73 (.I0(n2699), .I1(n2694), .I2(n2702), .I3(n2693), 
            .O(n37_c));
    defparam i14_4_lut_adj_73.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_74 (.I0(n2700), .I1(n36_adj_1866), .I2(n2687), 
            .I3(n2691), .O(n41_c));
    defparam i18_4_lut_adj_74.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n2698), .I1(n40_c), .I2(n32_adj_1867), .I3(n2692), 
            .O(n43_adj_1869));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43_adj_1869), .I1(n41_c), .I2(n37_c), .I3(n38_adj_1868), 
            .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20520_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25188));
    defparam i20520_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_155_add_1540_3_lut (.I0(n2212), .I1(n2212), .I2(n2225), 
            .I3(n22587), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_3_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i1004_1005 (.Q(n1191), .C(clock_c), .D(n11855));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1001_1002 (.Q(n1192), .C(clock_c), .D(n11854));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1004_11_lut (.I0(n1404_c), .I1(n1404_c), .I2(n1433_c), 
            .I3(n22463), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_17 (.CI(n22228), .I0(\ootx_payloads_N_1699[15] ), .I1(GND_net), 
            .CO(n22229));
    SB_CARRY add_154_13 (.CI(n22254), .I0(n2849[11]), .I1(GND_net), .CO(n22255));
    SB_CARRY mod_155_add_2076_28 (.CI(n22808), .I0(n2987), .I1(n3017), 
            .CO(n22809));
    SB_LUT4 mod_155_add_2009_24_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n22776), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_13_i1_3_lut (.I0(bit_counters_0_23), .I1(bit_counters_1_23), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[23]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_13_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i998_999 (.Q(n1193), .C(clock_c), .D(n11853));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i518_519 (.Q(ootx_payloads_0_80), .C(clock_c), .D(n11101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_adj_75 (.I0(n1108), .I1(n1103), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_1870));
    defparam i1_2_lut_adj_75.LUT_INIT = 16'heeee;
    SB_DFF i995_996 (.Q(n1194), .C(clock_c), .D(n11852));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i5_4_lut_adj_76 (.I0(n1106), .I1(n1107), .I2(n1104), .I3(n1105), 
            .O(n12));
    defparam i5_4_lut_adj_76.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_77 (.I0(n2851[21]), .I1(n1112), .I2(n1111), .I3(n1110), 
            .O(n22906));
    defparam i3_4_lut_adj_77.LUT_INIT = 16'hfffe;
    SB_DFF i992_993 (.Q(n1195), .C(clock_c), .D(n11851));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i989_990 (.Q(n1196), .C(clock_c), .D(n11850));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7562_3_lut_4_lut (.I0(n640), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1374), .O(n11672));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7562_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i986_987 (.Q(n1197), .C(clock_c), .D(n11849));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_2076_27_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n22807), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2076_27 (.CI(n22807), .I0(n2988), .I1(n3017), 
            .CO(n22808));
    SB_LUT4 i6970_3_lut_4_lut (.I0(n640), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_59), .O(n11080));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7012_3_lut_4_lut (.I0(n724), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_101), .O(n11122));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7012_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i983_984 (.Q(n1198), .C(clock_c), .D(n11848));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 PrioSelect_137_i2_3_lut (.I0(data), .I1(n4485[13]), .I2(n34[1]), 
            .I3(GND_net), .O(n170));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_137_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i980_981 (.Q(n1199), .C(clock_c), .D(n11847));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i977_978 (.Q(n1200), .C(clock_c), .D(n11846));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i974_975 (.Q(n1201), .C(clock_c), .D(n11845));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7706_3_lut_4_lut (.I0(n928), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1230), .O(n11816));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7706_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2009_24 (.CI(n22776), .I0(n2891), .I1(n2918), 
            .CO(n22777));
    SB_LUT4 mod_155_add_2009_23_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n22775), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i971_972 (.Q(n1202), .C(clock_c), .D(n11844));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i968_969 (.Q(n1203), .C(clock_c), .D(n11843));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i515_516 (.Q(ootx_payloads_0_79), .C(clock_c), .D(n11100));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i965_966 (.Q(n1204), .C(clock_c), .D(n11842));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2009_23 (.CI(n22775), .I0(n2892), .I1(n2918), 
            .CO(n22776));
    SB_LUT4 PrioSelect_133_i2_3_lut (.I0(data), .I1(n4485[12]), .I2(n34[1]), 
            .I3(GND_net), .O(n166));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_133_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i962_963 (.Q(n1205), .C(clock_c), .D(n11841));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1942_18 (.CI(n22743), .I0(n2797), .I1(n2819), 
            .CO(n22744));
    SB_LUT4 mod_155_add_1942_17_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n22742), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i959_960 (.Q(n1206), .C(clock_c), .D(n11840));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i956_957 (.Q(n1207), .C(clock_c), .D(n11839));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i953_954 (.Q(n1208), .C(clock_c), .D(n11838));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i6_4_lut (.I0(n22906), .I1(n12), .I2(n8_adj_1870), .I3(n1109), 
            .O(n1136));
    defparam i6_4_lut.LUT_INIT = 16'hfefc;
    SB_DFF i950_951 (.Q(n1209), .C(clock_c), .D(n11837));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i947_948 (.Q(n1210), .C(clock_c), .D(n11836));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7604_3_lut_4_lut (.I0(n724), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1332), .O(n11714));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7604_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1808_12_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n22686), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20521_1_lut (.I0(n1235_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25189));
    defparam i20521_1_lut.LUT_INIT = 16'h5555;
    SB_DFF i944_945 (.Q(n1211), .C(clock_c), .D(n11835));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i941_942 (.Q(n1212), .C(clock_c), .D(n11834));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7114_3_lut_4_lut (.I0(n928), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_203), .O(n11224));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7114_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i938_939 (.Q(n1213), .C(clock_c), .D(n11833));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1942_17 (.CI(n22742), .I0(n2798), .I1(n2819), 
            .CO(n22743));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_78 (.I0(n113), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n1010));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_78.LUT_INIT = 16'h0080;
    SB_DFF i935_936 (.Q(n1214), .C(clock_c), .D(n11832));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_79 (.I0(n113), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n754));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_79.LUT_INIT = 16'h0008;
    SB_LUT4 i7032_3_lut_4_lut (.I0(n764), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_121), .O(n11142));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7032_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1540_3 (.CI(n22587), .I0(n2212), .I1(n2225), 
            .CO(n22588));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_80 (.I0(n96), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n928));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_80.LUT_INIT = 16'h0080;
    SB_CARRY mod_155_add_1808_12 (.CI(n22686), .I0(n2603), .I1(n2621), 
            .CO(n22687));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_81 (.I0(n96), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n672));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_81.LUT_INIT = 16'h0008;
    SB_LUT4 PrioSelect_129_i2_3_lut (.I0(data), .I1(n4485[11]), .I2(n34[1]), 
            .I3(GND_net), .O(n162));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_129_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER ootx_states_0__i0_i1 (.Q(\ootx_states[0] [1]), .C(clock_c), 
            .E(n23163), .D(ootx_states_0__1__N_898[1]), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i7561_3_lut_4_lut (.I0(n638), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1375), .O(n11671));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_12_i1_3_lut (.I0(ootx_payloads_0_263), .I1(ootx_payloads_1_263), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[263]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 PrioSelect_125_i2_3_lut (.I0(data), .I1(n4485[10]), .I2(n34[1]), 
            .I3(GND_net), .O(n158));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_125_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6969_3_lut_4_lut (.I0(n638), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_58), .O(n11079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6969_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7705_3_lut_4_lut (.I0(n926), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1231), .O(n11815));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7705_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7113_3_lut_4_lut (.I0(n926), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_202), .O(n11223));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7113_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_82 (.I0(n94_adj_1872), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n926));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_82.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_83 (.I0(n94_adj_1872), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n670));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_83.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut_4_lut (.I0(n17_adj_1864), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n82_adj_1873));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i82_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i6256_4_lut (.I0(\lighthouse[0] ), .I1(ootx_payloads_N_1685), 
            .I2(n432), .I3(n17_c), .O(n10357));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i6256_4_lut.LUT_INIT = 16'h888a;
    SB_LUT4 i7624_3_lut_4_lut (.I0(n764), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1312), .O(n11734));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7624_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_84 (.I0(\lighthouse[0] ), .I1(n23_adj_1874), .I2(GND_net), 
            .I3(GND_net), .O(n20));
    defparam i1_2_lut_adj_84.LUT_INIT = 16'hdddd;
    SB_LUT4 Mux_13_i1_3_lut_adj_85 (.I0(ootx_payloads_0_262), .I1(ootx_payloads_1_262), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[262]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_13_i1_3_lut_adj_85.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut_4_lut (.I0(n17_adj_1864), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n81));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i81_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i7704_3_lut_4_lut (.I0(n924), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1232), .O(n11814));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7704_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7112_3_lut_4_lut (.I0(n924), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_201), .O(n11222));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7112_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7560_3_lut_4_lut (.I0(n636), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1376), .O(n11670));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6968_3_lut_4_lut (.I0(n636), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_57), .O(n11078));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6968_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_86 (.I0(n92), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n924));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_86.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_87 (.I0(n92), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n668));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_87.LUT_INIT = 16'h0008;
    SB_LUT4 i7703_3_lut_4_lut (.I0(n922), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1233), .O(n11813));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7703_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7111_3_lut_4_lut (.I0(n922), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_200), .O(n11221));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7111_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7559_3_lut_4_lut (.I0(n634), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1377), .O(n11669));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7559_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6967_3_lut_4_lut (.I0(n634), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_56), .O(n11077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6967_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_88 (.I0(n90_adj_1876), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n922));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_88.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_89 (.I0(n90_adj_1876), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n666));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_89.LUT_INIT = 16'h0008;
    SB_LUT4 i7702_3_lut_4_lut (.I0(n920), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1234), .O(n11812));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7702_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7110_3_lut_4_lut (.I0(n920), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_199), .O(n11220));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7110_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7558_3_lut_4_lut (.I0(n632), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1378), .O(n11668));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6966_3_lut_4_lut (.I0(n632), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_55), .O(n11076));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6966_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_90 (.I0(n88_adj_1877), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n920));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_90.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_91 (.I0(n88_adj_1877), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n664));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_91.LUT_INIT = 16'h0008;
    SB_LUT4 i7701_3_lut_4_lut (.I0(n918), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1235), .O(n11811));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7701_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7109_3_lut_4_lut (.I0(n918), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_198), .O(n11219));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7109_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_92 (.I0(n86_adj_1860), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n918));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_92.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_93 (.I0(n86_adj_1860), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n662));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_93.LUT_INIT = 16'h0008;
    SB_LUT4 i7700_3_lut_4_lut (.I0(n916), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1236), .O(n11810));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7700_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7108_3_lut_4_lut (.I0(n916), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_197), .O(n11218));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7108_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7026_3_lut_4_lut (.I0(n752), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_115), .O(n11136));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7026_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7618_3_lut_4_lut (.I0(n752), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1318), .O(n11728));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7618_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_94 (.I0(n84), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n916));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_94.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_95 (.I0(n84), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n660));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_95.LUT_INIT = 16'h0008;
    SB_LUT4 i7699_3_lut_4_lut (.I0(n914), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1237), .O(n11809));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7699_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7107_3_lut_4_lut (.I0(n914), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_196), .O(n11217));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7107_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_96 (.I0(n82_adj_1873), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n914));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_96.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_97 (.I0(n82_adj_1873), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n658));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_97.LUT_INIT = 16'h0008;
    SB_LUT4 i2_3_lut_adj_98 (.I0(ootx_payloads_N_1744[0]), .I1(new_data), 
            .I2(ootx_payloads_N_1744[1]), .I3(GND_net), .O(n4729));
    defparam i2_3_lut_adj_98.LUT_INIT = 16'h0404;
    SB_LUT4 i7581_3_lut_4_lut (.I0(n678), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1355), .O(n11691));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7581_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_99 (.I0(reset_c), .I1(n4729), .I2(GND_net), .I3(GND_net), 
            .O(ootx_shift_registers_N_1748));
    defparam i1_2_lut_adj_99.LUT_INIT = 16'h4444;
    SB_LUT4 i7698_3_lut_4_lut (.I0(n912), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1238), .O(n11808));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7698_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7106_3_lut_4_lut (.I0(n912), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_195), .O(n11216));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7106_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_365_i1_3_lut (.I0(ootx_shift_registers_0_13), .I1(ootx_shift_registers_1_13), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[13]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_365_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_378_i1_3_lut (.I0(ootx_shift_registers_0_0), .I1(ootx_shift_registers_1_0), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_378_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_364_i1_3_lut (.I0(ootx_shift_registers_0_14), .I1(ootx_shift_registers_1_14), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[14]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_364_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_372_i1_3_lut (.I0(ootx_shift_registers_0_6), .I1(ootx_shift_registers_1_6), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[6]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_372_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_369_i1_3_lut (.I0(ootx_shift_registers_0_9), .I1(ootx_shift_registers_1_9), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[9]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_369_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_363_i1_3_lut (.I0(ootx_shift_registers_0_15), .I1(ootx_shift_registers_1_15), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[15]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_363_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(ootx_shift_registers_0_10), .I1(data_counters_N_1780[13]), 
            .I2(ootx_shift_registers_1_10), .I3(\lighthouse[0] ), .O(n20_adj_1881));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i2_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 Mux_374_i1_3_lut (.I0(ootx_shift_registers_0_4), .I1(ootx_shift_registers_1_4), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[4]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_374_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_100 (.I0(ootx_shift_registers_0_2), .I1(data_counters_N_1780[15]), 
            .I2(ootx_shift_registers_1_2), .I3(\lighthouse[0] ), .O(n19_adj_1882));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i1_4_lut_adj_100.LUT_INIT = 16'hfcee;
    SB_LUT4 Mux_361_i1_3_lut (.I0(ootx_shift_registers_0_17), .I1(ootx_shift_registers_1_17), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[17]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_361_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_371_i1_3_lut (.I0(ootx_shift_registers_0_7), .I1(ootx_shift_registers_1_7), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[7]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_371_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_362_i1_3_lut (.I0(ootx_shift_registers_0_16), .I1(ootx_shift_registers_1_16), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(data_counters_N_1780[16]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[31:41])
    defparam Mux_362_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_101 (.I0(ootx_shift_registers_0_11), .I1(data_counters_N_1780[0]), 
            .I2(ootx_shift_registers_1_11), .I3(\lighthouse[0] ), .O(n24_adj_1883));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i6_4_lut_adj_101.LUT_INIT = 16'hf3bb;
    SB_LUT4 i4_4_lut_adj_102 (.I0(ootx_shift_registers_0_12), .I1(data_counters_N_1780[14]), 
            .I2(ootx_shift_registers_1_12), .I3(\lighthouse[0] ), .O(n22_adj_1884));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i4_4_lut_adj_102.LUT_INIT = 16'hfcee;
    SB_LUT4 i5_4_lut_adj_103 (.I0(ootx_shift_registers_0_5), .I1(data_counters_N_1780[6]), 
            .I2(ootx_shift_registers_1_5), .I3(\lighthouse[0] ), .O(n23_adj_1885));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i5_4_lut_adj_103.LUT_INIT = 16'hfcee;
    SB_LUT4 i7557_3_lut_4_lut (.I0(n630), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1379), .O(n11667));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_14_i1_3_lut_adj_104 (.I0(ootx_payloads_0_261), .I1(ootx_payloads_1_261), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[261]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_14_i1_3_lut_adj_104.LUT_INIT = 16'hcaca;
    SB_LUT4 i6965_3_lut_4_lut (.I0(n630), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_54), .O(n11075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6965_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_15_i1_3_lut_adj_105 (.I0(ootx_payloads_0_260), .I1(ootx_payloads_1_260), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[260]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_15_i1_3_lut_adj_105.LUT_INIT = 16'hcaca;
    SB_LUT4 i6989_3_lut_4_lut (.I0(n678), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_78), .O(n11099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 PrioSelect_121_i2_3_lut (.I0(data), .I1(n4485[9]), .I2(n34[1]), 
            .I3(GND_net), .O(n154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_121_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_106 (.I0(n80), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n912));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_106.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_107 (.I0(n80), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n656));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_107.LUT_INIT = 16'h0008;
    SB_LUT4 Mux_16_i1_3_lut_adj_108 (.I0(ootx_payloads_0_259), .I1(ootx_payloads_1_259), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[259]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_16_i1_3_lut_adj_108.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_2076_26_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n22806), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7697_3_lut_4_lut (.I0(n910), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1239), .O(n11807));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7697_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_109 (.I0(ootx_shift_registers_0_1), .I1(data_counters_N_1780[16]), 
            .I2(ootx_shift_registers_1_1), .I3(\lighthouse[0] ), .O(n21));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i3_4_lut_adj_109.LUT_INIT = 16'hfcee;
    SB_LUT4 i8_4_lut_adj_110 (.I0(ootx_shift_registers_0_3), .I1(data_counters_N_1780[9]), 
            .I2(ootx_shift_registers_1_3), .I3(\lighthouse[0] ), .O(n26_adj_1887));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i8_4_lut_adj_110.LUT_INIT = 16'hfcee;
    SB_LUT4 i14_4_lut_adj_111 (.I0(data_counters_N_1780[17]), .I1(n19_adj_1882), 
            .I2(data_counters_N_1780[4]), .I3(n20_adj_1881), .O(n32_adj_1888));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i14_4_lut_adj_111.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_112 (.I0(ootx_shift_registers_0_8), .I1(data_counters_N_1780[7]), 
            .I2(ootx_shift_registers_1_8), .I3(\lighthouse[0] ), .O(n25_adj_1889));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i7_4_lut_adj_112.LUT_INIT = 16'hfcee;
    SB_LUT4 i15_4_lut_adj_113 (.I0(n21), .I1(n23_adj_1885), .I2(n22_adj_1884), 
            .I3(n24_adj_1883), .O(n33_adj_1890));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i15_4_lut_adj_113.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_114 (.I0(n33_adj_1890), .I1(n25_adj_1889), .I2(n32_adj_1888), 
            .I3(n26_adj_1887), .O(n35));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam i17_4_lut_adj_114.LUT_INIT = 16'hfffe;
    SB_LUT4 i7105_3_lut_4_lut (.I0(n910), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_194), .O(n11215));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7105_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19466_3_lut (.I0(crc32s_N_1751), .I1(n432), .I2(ootx_payloads_N_1685), 
            .I3(GND_net), .O(n24133));
    defparam i19466_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_115 (.I0(n17_c), .I1(n1119), .I2(n24133), .I3(data_counters_N_1776), 
            .O(n23_adj_1874));
    defparam i1_4_lut_adj_115.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_116 (.I0(ootx_payloads_N_1744[1]), .I1(ootx_payloads_N_1744[0]), 
            .I2(GND_net), .I3(GND_net), .O(n118));
    defparam i1_2_lut_adj_116.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_117 (.I0(ootx_payloads_N_1699[2]), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(ootx_payloads_N_1699[1]), .I3(GND_net), .O(n8941));
    defparam i2_3_lut_adj_117.LUT_INIT = 16'h8080;
    SB_LUT4 Mux_22_i1_3_lut (.I0(data_counters_0_16), .I1(data_counters_1_16), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[16]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_15_i1_3_lut_adj_118 (.I0(data_counters_0_23), .I1(data_counters_1_23), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[23]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_15_i1_3_lut_adj_118.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_10_i1_3_lut (.I0(data_counters_0_28), .I1(data_counters_1_28), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[28]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_10_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_18_i1_3_lut_adj_119 (.I0(data_counters_0_20), .I1(data_counters_1_20), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[20]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_18_i1_3_lut_adj_119.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_120 (.I0(n78_adj_1891), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n910));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_120.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_121 (.I0(n78_adj_1891), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n654));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_121.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_122 (.I0(n111), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n1008));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_122.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_123 (.I0(n111), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n752));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_123.LUT_INIT = 16'h0008;
    SB_LUT4 i7580_3_lut_4_lut (.I0(n676), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1356), .O(n11690));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7580_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7696_3_lut_4_lut (.I0(n908), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1240), .O(n11806));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7696_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_17_i1_3_lut_adj_124 (.I0(ootx_payloads_0_258), .I1(ootx_payloads_1_258), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[258]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_17_i1_3_lut_adj_124.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_2009_22_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n22774), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7104_3_lut_4_lut (.I0(n908), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_193), .O(n11214));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7104_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2076_26 (.CI(n22806), .I0(n2989), .I1(n3017), 
            .CO(n22807));
    SB_LUT4 Mux_18_i1_3_lut_adj_125 (.I0(ootx_payloads_0_257), .I1(ootx_payloads_1_257), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[257]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_18_i1_3_lut_adj_125.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_19_i1_3_lut_adj_126 (.I0(ootx_payloads_0_256), .I1(ootx_payloads_1_256), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[256]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_19_i1_3_lut_adj_126.LUT_INIT = 16'hcaca;
    SB_LUT4 i7556_3_lut_4_lut (.I0(n628), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1380), .O(n11666));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7556_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_20_i1_3_lut (.I0(ootx_payloads_0_255), .I1(ootx_payloads_1_255), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[255]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_20_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2009_22 (.CI(n22774), .I0(n2893), .I1(n2918), 
            .CO(n22775));
    SB_LUT4 PrioSelect_117_i2_3_lut (.I0(data), .I1(n4485[8]), .I2(n34[1]), 
            .I3(GND_net), .O(n150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_117_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_19_i1_3_lut_adj_127 (.I0(data_counters_0_19), .I1(data_counters_1_19), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[19]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_19_i1_3_lut_adj_127.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_16_i1_3_lut_adj_128 (.I0(data_counters_0_22), .I1(data_counters_1_22), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[22]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_16_i1_3_lut_adj_128.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_11_i1_3_lut (.I0(data_counters_0_27), .I1(data_counters_1_27), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[27]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_11_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_17_i1_3_lut_adj_129 (.I0(data_counters_0_21), .I1(data_counters_1_21), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[21]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_17_i1_3_lut_adj_129.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_13_i1_3_lut_adj_130 (.I0(data_counters_0_25), .I1(data_counters_1_25), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[25]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_13_i1_3_lut_adj_130.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_12_i1_3_lut_adj_131 (.I0(data_counters_0_26), .I1(data_counters_1_26), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[26]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_12_i1_3_lut_adj_131.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_9_i1_3_lut (.I0(data_counters_0_29), .I1(data_counters_1_29), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[29]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_9_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_14_i1_3_lut_adj_132 (.I0(data_counters_0_24), .I1(data_counters_1_24), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[24]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_14_i1_3_lut_adj_132.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_8_i1_3_lut (.I0(data_counters_0_30), .I1(data_counters_1_30), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[30] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_8_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_133 (.I0(ootx_payloads_N_1699[28]), .I1(ootx_payloads_N_1699[23]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_1895));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i1_2_lut_adj_133.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_134 (.I0(ootx_payloads_N_1699[24]), .I1(ootx_payloads_N_1699[29]), 
            .I2(ootx_payloads_N_1699[26]), .I3(n10_adj_1895), .O(n16_adj_1896));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i7_4_lut_adj_134.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_135 (.I0(ootx_payloads_N_1699[25]), .I1(ootx_payloads_N_1699[21]), 
            .I2(ootx_payloads_N_1699[27]), .I3(ootx_payloads_N_1699[22]), 
            .O(n15));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i6_4_lut_adj_135.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_136 (.I0(n15), .I1(ootx_payloads_N_1699[19]), .I2(n16_adj_1896), 
            .I3(ootx_payloads_N_1699[20]), .O(n4_adj_1897));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i1_4_lut_adj_136.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_137 (.I0(ootx_payloads_N_1699[17]), .I1(n4_adj_1897), 
            .I2(ootx_payloads_N_1699[16]), .I3(ootx_payloads_N_1699[18]), 
            .O(n9200));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i2_4_lut_adj_137.LUT_INIT = 16'hfffe;
    SB_LUT4 Mux_29_i1_3_lut_adj_138 (.I0(data_counters_0_9), .I1(data_counters_1_9), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[9] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_29_i1_3_lut_adj_138.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_25_i1_3_lut (.I0(data_counters_0_13), .I1(data_counters_1_13), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[13] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_25_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_26_i1_3_lut_adj_139 (.I0(data_counters_0_12), .I1(data_counters_1_12), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[12] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_26_i1_3_lut_adj_139.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_27_i1_3_lut_adj_140 (.I0(data_counters_0_11), .I1(data_counters_1_11), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[11] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_27_i1_3_lut_adj_140.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_21_i1_3_lut (.I0(ootx_payloads_0_254), .I1(ootx_payloads_1_254), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[254]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6964_3_lut_4_lut (.I0(n628), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_53), .O(n11074));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6964_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_22_i1_3_lut_adj_141 (.I0(ootx_payloads_0_253), .I1(ootx_payloads_1_253), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[253]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_22_i1_3_lut_adj_141.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_142 (.I0(n76), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n908));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_142.LUT_INIT = 16'h0080;
    SB_LUT4 Mux_23_i1_3_lut (.I0(ootx_payloads_0_252), .I1(ootx_payloads_1_252), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[252]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_23_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_143 (.I0(\lighthouse[0] ), .I1(n4729), .I2(GND_net), 
            .I3(GND_net), .O(n23741));
    defparam i1_2_lut_adj_143.LUT_INIT = 16'h8888;
    SB_LUT4 i6988_3_lut_4_lut (.I0(n676), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_77), .O(n11098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6988_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_24_i1_3_lut (.I0(ootx_payloads_0_251), .I1(ootx_payloads_1_251), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[251]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_24_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_144 (.I0(n76), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n652));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_144.LUT_INIT = 16'h0008;
    SB_LUT4 i7695_3_lut_4_lut (.I0(n906), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1241), .O(n11805));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7695_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_25_i1_3_lut_adj_145 (.I0(ootx_payloads_0_250), .I1(ootx_payloads_1_250), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[250]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_25_i1_3_lut_adj_145.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_26_i1_3_lut_adj_146 (.I0(ootx_payloads_0_249), .I1(ootx_payloads_1_249), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[249]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_26_i1_3_lut_adj_146.LUT_INIT = 16'hcaca;
    SB_LUT4 i7103_3_lut_4_lut (.I0(n906), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_192), .O(n11213));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7103_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_147 (.I0(n74_adj_1899), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n906));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_147.LUT_INIT = 16'h0080;
    SB_LUT4 Mux_28_i1_3_lut_adj_148 (.I0(data_counters_0_10), .I1(data_counters_1_10), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[10] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_28_i1_3_lut_adj_148.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_24_i1_3_lut_adj_149 (.I0(data_counters_0_14), .I1(data_counters_1_14), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[14] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_24_i1_3_lut_adj_149.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(\ootx_payloads_N_1699[15] ), .I1(\ootx_payloads_N_1699[14] ), 
            .I2(\ootx_payloads_N_1699[10] ), .I3(GND_net), .O(n14));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_2_lut (.I0(\ootx_payloads_N_1699[11] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_1900));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_150 (.I0(\ootx_payloads_N_1699[12] ), .I1(\ootx_payloads_N_1699[8] ), 
            .I2(\ootx_payloads_N_1699[13] ), .I3(\ootx_payloads_N_1699[9] ), 
            .O(n15_adj_1901));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(118[10:40])
    defparam i6_4_lut_adj_150.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_151 (.I0(\ootx_payloads_N_1699[6] ), .I1(n15_adj_1901), 
            .I2(n13_adj_1900), .I3(n14), .O(n24013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[11:42])
    defparam i1_4_lut_adj_151.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_152 (.I0(\ootx_payloads_N_1699[5] ), .I1(n9200), 
            .I2(\ootx_payloads_N_1699[30] ), .I3(n24013), .O(n24018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_4_lut_adj_152.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_153 (.I0(n74_adj_1899), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n650));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_153.LUT_INIT = 16'h0008;
    SB_LUT4 i7555_3_lut_4_lut (.I0(n626), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1381), .O(n11665));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7555_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6963_3_lut_4_lut (.I0(n626), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_52), .O(n11073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6963_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7694_3_lut_4_lut (.I0(n904), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1242), .O(n11804));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7694_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7102_3_lut_4_lut (.I0(n904), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_191), .O(n11212));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7102_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i135_2_lut_3_lut (.I0(n39_adj_1902), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n135));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i135_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut_4_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n80));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i80_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut_4_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n79));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i79_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_154 (.I0(n135), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n904));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_154.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_155 (.I0(n135), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n648));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_155.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i136_2_lut_3_lut (.I0(n39_adj_1902), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n136));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i136_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 PrioSelect_113_i2_3_lut (.I0(data), .I1(n4485[7]), .I2(n34[1]), 
            .I3(GND_net), .O(n146));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_113_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7732_3_lut_4_lut (.I0(n980), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1204), .O(n11842));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7732_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7554_3_lut_4_lut (.I0(n624), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1382), .O(n11664));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7554_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_27_i1_3_lut_adj_156 (.I0(ootx_payloads_0_248), .I1(ootx_payloads_1_248), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[248]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_27_i1_3_lut_adj_156.LUT_INIT = 16'hcaca;
    SB_LUT4 i7140_3_lut_4_lut (.I0(n980), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_229), .O(n11250));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7140_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6962_3_lut_4_lut (.I0(n624), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_51), .O(n11072));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6962_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 PrioSelect_109_i2_3_lut (.I0(data), .I1(n4485[6]), .I2(n34[1]), 
            .I3(GND_net), .O(n142));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_109_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_28_i1_3_lut_adj_157 (.I0(ootx_payloads_0_247), .I1(ootx_payloads_1_247), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[247]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_28_i1_3_lut_adj_157.LUT_INIT = 16'hcaca;
    SB_LUT4 i7693_3_lut_4_lut (.I0(n902), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1243), .O(n11803));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7693_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut (.I0(n20112), .I1(n23985), .I2(n20105), .I3(GND_net), 
            .O(n432));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i1_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i1_2_lut_adj_158 (.I0(new_data), .I1(reset_c), .I2(GND_net), 
            .I3(GND_net), .O(n9498));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_adj_158.LUT_INIT = 16'h2222;
    SB_LUT4 i7101_3_lut_4_lut (.I0(n902), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_190), .O(n11211));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7101_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7692_3_lut_4_lut (.I0(n900), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1244), .O(n11802));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7692_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7100_3_lut_4_lut (.I0(n900), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_189), .O(n11210));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7100_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6126_4_lut (.I0(\lighthouse[0] ), .I1(ootx_payloads_N_1685), 
            .I2(n432), .I3(n17_c), .O(n10243));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(54[9:22])
    defparam i6126_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 EnabledDecoder_2_i162_2_lut_3_lut (.I0(n66_adj_1904), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n162_adj_1905));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i162_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i7731_3_lut_4_lut (.I0(n978), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1205), .O(n11841));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7731_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7139_3_lut_4_lut (.I0(n978), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_228), .O(n11249));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7139_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7579_3_lut_4_lut (.I0(n674), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1357), .O(n11689));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7579_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_159 (.I0(\lighthouse[0] ), .I1(n23_adj_1874), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i1_2_lut_adj_159.LUT_INIT = 16'heeee;
    SB_LUT4 i7553_3_lut_4_lut (.I0(n622), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1383), .O(n11663));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7553_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_29_i1_3_lut_adj_160 (.I0(ootx_payloads_0_246), .I1(ootx_payloads_1_246), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[246]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_29_i1_3_lut_adj_160.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_30_i1_3_lut (.I0(ootx_payloads_0_245), .I1(ootx_payloads_1_245), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[245]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_30_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6961_3_lut_4_lut (.I0(n622), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_50), .O(n11071));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6961_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7691_3_lut_4_lut (.I0(n898), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1245), .O(n11801));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7691_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_31_i1_3_lut (.I0(ootx_payloads_0_244), .I1(ootx_payloads_1_244), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[244]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_31_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7099_3_lut_4_lut (.I0(n898), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_188), .O(n11209));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7099_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7690_3_lut_4_lut (.I0(n896), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1246), .O(n11800));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7690_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7098_3_lut_4_lut (.I0(n896), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_187), .O(n11208));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7098_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1004_11 (.CI(n22463), .I0(n1404_c), .I1(n1433_c), 
            .CO(n22464));
    SB_CARRY add_355_13 (.CI(n22285), .I0(\counter_from_last_rise[11] ), 
            .I1(GND_net), .CO(n22286));
    SB_LUT4 mod_155_add_1540_2_lut (.I0(n2851[10]), .I1(n2851[10]), .I2(n25179), 
            .I3(VCC_net), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i7552_3_lut_4_lut (.I0(n620), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1384), .O(n11662));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_355_12_lut (.I0(GND_net), .I1(\counter_from_last_rise[10] ), 
            .I2(GND_net), .I3(n22284), .O(n6355)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6960_3_lut_4_lut (.I0(n620), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_49), .O(n11070));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6960_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7689_3_lut_4_lut (.I0(n894), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1247), .O(n11799));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7689_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7097_3_lut_4_lut (.I0(n894), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_186), .O(n11207));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7097_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1808_11_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n22685), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1004_10_lut (.I0(n1405_c), .I1(n1405_c), .I2(n1433_c), 
            .I3(n22462), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_12 (.CI(n22284), .I0(\counter_from_last_rise[10] ), 
            .I1(GND_net), .CO(n22285));
    SB_LUT4 add_355_11_lut (.I0(GND_net), .I1(\counter_from_last_rise[9] ), 
            .I2(GND_net), .I3(n22283), .O(n6356)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1808_11 (.CI(n22685), .I0(n2604), .I1(n2621), 
            .CO(n22686));
    SB_LUT4 mod_155_add_1942_16_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n22741), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_10_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n22684), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1540_2 (.CI(VCC_net), .I0(n2851[10]), .I1(n25179), 
            .CO(n22587));
    SB_CARRY add_355_11 (.CI(n22283), .I0(\counter_from_last_rise[9] ), 
            .I1(GND_net), .CO(n22284));
    SB_LUT4 add_154_12_lut (.I0(GND_net), .I1(n2849[10]), .I2(GND_net), 
            .I3(n22253), .O(n2851[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1004_10 (.CI(n22462), .I0(n1405_c), .I1(n1433_c), 
            .CO(n22463));
    SB_CARRY add_154_12 (.CI(n22253), .I0(n2849[10]), .I1(GND_net), .CO(n22254));
    SB_LUT4 add_355_10_lut (.I0(GND_net), .I1(\counter_from_last_rise[8] ), 
            .I2(GND_net), .I3(n22282), .O(n6357)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_161 (.I0(n125), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n894));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_161.LUT_INIT = 16'h0020;
    SB_LUT4 mod_155_add_1473_22_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n22586), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_11_lut (.I0(GND_net), .I1(n2849[9]), .I2(GND_net), 
            .I3(n22252), .O(n2851[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_66_16_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[14] ), 
            .I2(GND_net), .I3(n22227), .O(n337[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1004_9_lut (.I0(n1406_c), .I1(n1406_c), .I2(n1433_c), 
            .I3(n22461), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_5 (.CI(n22216), .I0(\ootx_payloads_N_1699[3] ), .I1(GND_net), 
            .CO(n22217));
    SB_LUT4 Mux_16_i1_3_lut_adj_162 (.I0(payload_lengths_0_4), .I1(payload_lengths_1_4), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[4] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_16_i1_3_lut_adj_162.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_163 (.I0(n125), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n638));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_163.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_1942_16 (.CI(n22741), .I0(n2799), .I1(n2819), 
            .CO(n22742));
    SB_CARRY add_66_16 (.CI(n22227), .I0(\ootx_payloads_N_1699[14] ), .I1(GND_net), 
            .CO(n22228));
    SB_CARRY add_154_11 (.CI(n22252), .I0(n2849[9]), .I1(GND_net), .CO(n22253));
    SB_CARRY mod_155_add_1808_10 (.CI(n22684), .I0(n2605), .I1(n2621), 
            .CO(n22685));
    SB_LUT4 mod_155_add_1808_9_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n22683), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_10 (.CI(n22282), .I0(\counter_from_last_rise[8] ), 
            .I1(GND_net), .CO(n22283));
    SB_LUT4 mod_155_add_2076_25_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n22805), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_21_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n22585), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_10_lut (.I0(GND_net), .I1(n2849[8]), .I2(GND_net), 
            .I3(n22251), .O(n2851[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_154_10 (.CI(n22251), .I0(n2849[8]), .I1(GND_net), .CO(n22252));
    SB_CARRY mod_155_add_1004_9 (.CI(n22461), .I0(n1406_c), .I1(n1433_c), 
            .CO(n22462));
    SB_LUT4 add_355_9_lut (.I0(GND_net), .I1(\counter_from_last_rise[7] ), 
            .I2(GND_net), .I3(n22281), .O(n6358)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_154_9_lut (.I0(GND_net), .I1(n2849[7]), .I2(GND_net), 
            .I3(n22250), .O(n2851[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7025_3_lut_4_lut (.I0(n750), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_114), .O(n11135));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7617_3_lut_4_lut (.I0(n750), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1319), .O(n11727));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7617_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1473_21 (.CI(n22585), .I0(n2094), .I1(n2126), 
            .CO(n22586));
    SB_LUT4 add_66_15_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[13] ), 
            .I2(GND_net), .I3(n22226), .O(n337[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7551_3_lut_4_lut (.I0(n618), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1385), .O(n11661));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6959_3_lut_4_lut (.I0(n618), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_48), .O(n11069));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6959_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7688_3_lut_4_lut (.I0(n892), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1248), .O(n11798));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7688_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1004_8_lut (.I0(n1407_c), .I1(n1407_c), .I2(n1433_c), 
            .I3(n22460), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_15 (.CI(n22226), .I0(\ootx_payloads_N_1699[13] ), .I1(GND_net), 
            .CO(n22227));
    SB_CARRY mod_155_add_1808_9 (.CI(n22683), .I0(n2606), .I1(n2621), 
            .CO(n22684));
    SB_CARRY add_154_9 (.CI(n22250), .I0(n2849[7]), .I1(GND_net), .CO(n22251));
    SB_LUT4 mod_155_add_2009_21_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n22773), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_20_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n22584), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_15_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n22740), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_8_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n22682), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7096_3_lut_4_lut (.I0(n892), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_185), .O(n11206));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7096_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_164 (.I0(\lighthouse[0] ), .I1(n23989), .I2(n4729), 
            .I3(n23985), .O(n23990));
    defparam i1_4_lut_adj_164.LUT_INIT = 16'hc8c0;
    SB_CARRY mod_155_add_1004_8 (.CI(n22460), .I0(n1407_c), .I1(n1433_c), 
            .CO(n22461));
    SB_CARRY add_355_9 (.CI(n22281), .I0(\counter_from_last_rise[7] ), .I1(GND_net), 
            .CO(n22282));
    SB_LUT4 add_355_8_lut (.I0(GND_net), .I1(\counter_from_last_rise[6] ), 
            .I2(GND_net), .I3(n22280), .O(n6359)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1473_20 (.CI(n22584), .I0(n2095), .I1(n2126), 
            .CO(n22585));
    SB_CARRY mod_155_add_1808_8 (.CI(n22682), .I0(n2607), .I1(n2621), 
            .CO(n22683));
    SB_CARRY add_355_8 (.CI(n22280), .I0(\counter_from_last_rise[6] ), .I1(GND_net), 
            .CO(n22281));
    SB_LUT4 mod_155_add_1004_7_lut (.I0(n1408_c), .I1(n1408_c), .I2(n1433_c), 
            .I3(n22459), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_355_7_lut (.I0(GND_net), .I1(counter_from_last_rise_c[5]), 
            .I2(GND_net), .I3(n22279), .O(n6333_c[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1942_15 (.CI(n22740), .I0(n2800), .I1(n2819), 
            .CO(n22741));
    SB_CARRY mod_155_add_2009_21 (.CI(n22773), .I0(n2894), .I1(n2918), 
            .CO(n22774));
    SB_LUT4 mod_155_add_1808_7_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n22681), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_7 (.CI(n22279), .I0(counter_from_last_rise_c[5]), .I1(GND_net), 
            .CO(n22280));
    SB_LUT4 Mux_32_i1_3_lut (.I0(ootx_payloads_0_243), .I1(ootx_payloads_1_243), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[243]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_32_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1942_14_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n22739), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_8_lut (.I0(GND_net), .I1(n2849[6]), .I2(GND_net), 
            .I3(n22249), .O(n2851[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_154_8 (.CI(n22249), .I0(n2849[6]), .I1(GND_net), .CO(n22250));
    SB_CARRY mod_155_add_1808_7 (.CI(n22681), .I0(n2608), .I1(n2621), 
            .CO(n22682));
    SB_LUT4 add_355_6_lut (.I0(GND_net), .I1(counter_from_last_rise[4]), 
            .I2(GND_net), .I3(n22278), .O(n6361)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_154_7_lut (.I0(GND_net), .I1(n2849[5]), .I2(GND_net), 
            .I3(n22248), .O(n2851[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1473_19_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n22583), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_14_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[12] ), 
            .I2(GND_net), .I3(n22225), .O(n337[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1004_7 (.CI(n22459), .I0(n1408_c), .I1(n1433_c), 
            .CO(n22460));
    SB_LUT4 i7687_3_lut_4_lut (.I0(n890), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1249), .O(n11797));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7687_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_33_i1_3_lut (.I0(ootx_payloads_0_242), .I1(ootx_payloads_1_242), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[242]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_33_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_165 (.I0(n2851[2]), .I1(n3012), .I2(n3011), .I3(n3010), 
            .O(n22903));
    defparam i3_4_lut_adj_165.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_166 (.I0(n22903), .I1(n2986), .I2(n3009), .I3(GND_net), 
            .O(n30_adj_1907));
    defparam i4_3_lut_adj_166.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_167 (.I0(n2999), .I1(n2990), .I2(n3005), .I3(n3006), 
            .O(n42_c));
    defparam i16_4_lut_adj_167.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_168 (.I0(n2996), .I1(n3000), .I2(n2987), .I3(n3001), 
            .O(n40_adj_1908));
    defparam i14_4_lut_adj_168.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_169 (.I0(n2994), .I1(n3003), .I2(n3004), .I3(n2992), 
            .O(n45_c));
    defparam i19_4_lut_adj_169.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_170 (.I0(n2984), .I1(n3007), .I2(n2991), .I3(n2993), 
            .O(n44_c));
    defparam i18_4_lut_adj_170.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_171 (.I0(n2985), .I1(n2995), .I2(n2997), .I3(n2998), 
            .O(n43_adj_1909));
    defparam i17_4_lut_adj_171.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n3002), .I1(n42_c), .I2(n30_adj_1907), .I3(n2988), 
            .O(n47_c));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1473_19 (.CI(n22583), .I0(n2096), .I1(n2126), 
            .CO(n22584));
    SB_CARRY add_66_14 (.CI(n22225), .I0(\ootx_payloads_N_1699[12] ), .I1(GND_net), 
            .CO(n22226));
    SB_CARRY add_154_7 (.CI(n22248), .I0(n2849[5]), .I1(GND_net), .CO(n22249));
    SB_LUT4 mod_155_add_1004_6_lut (.I0(n1409_c), .I1(n1409_c), .I2(n25184), 
            .I3(n22458), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1808_6_lut (.I0(n2609), .I1(n2609), .I2(n25178), 
            .I3(n22680), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_355_6 (.CI(n22278), .I0(counter_from_last_rise[4]), .I1(GND_net), 
            .CO(n22279));
    SB_LUT4 i7095_3_lut_4_lut (.I0(n890), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_184), .O(n11205));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7095_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1808_6 (.CI(n22680), .I0(n2609), .I1(n25178), 
            .CO(n22681));
    SB_LUT4 i6987_3_lut_4_lut (.I0(n674), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_76), .O(n11097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6987_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_154_6_lut (.I0(GND_net), .I1(n2849[4]), .I2(GND_net), 
            .I3(n22247), .O(n2851[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_154_6 (.CI(n22247), .I0(n2849[4]), .I1(GND_net), .CO(n22248));
    SB_LUT4 mod_155_add_1473_18_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n22582), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_355_5_lut (.I0(GND_net), .I1(counter_from_last_rise[3]), 
            .I2(GND_net), .I3(n22277), .O(n6362)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_154_5_lut (.I0(GND_net), .I1(n2849[3]), .I2(GND_net), 
            .I3(n22246), .O(n2851[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7550_3_lut_4_lut (.I0(n616), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1386), .O(n11660));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1004_6 (.CI(n22458), .I0(n1409_c), .I1(n25184), 
            .CO(n22459));
    SB_LUT4 add_66_13_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[11] ), 
            .I2(GND_net), .I3(n22224), .O(n337[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6958_3_lut_4_lut (.I0(n616), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_47), .O(n11068));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6958_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1473_18 (.CI(n22582), .I0(n2097), .I1(n2126), 
            .CO(n22583));
    SB_CARRY add_66_4 (.CI(n22215), .I0(ootx_payloads_N_1699[2]), .I1(GND_net), 
            .CO(n22216));
    SB_LUT4 i1_4_lut_adj_172 (.I0(n24110), .I1(n23989), .I2(n4729), .I3(n4), 
            .O(n23992));
    defparam i1_4_lut_adj_172.LUT_INIT = 16'hc4c0;
    SB_LUT4 mod_155_add_1004_5_lut (.I0(n1410_c), .I1(n1410_c), .I2(n1433_c), 
            .I3(n22457), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_13 (.CI(n22224), .I0(\ootx_payloads_N_1699[11] ), .I1(GND_net), 
            .CO(n22225));
    SB_CARRY add_154_5 (.CI(n22246), .I0(n2849[3]), .I1(GND_net), .CO(n22247));
    SB_CARRY mod_155_add_1942_14 (.CI(n22739), .I0(n2801), .I1(n2819), 
            .CO(n22740));
    SB_LUT4 mod_155_add_2143_33_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n22842), .O(n63_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_33_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2076_25 (.CI(n22805), .I0(n2990), .I1(n3017), 
            .CO(n22806));
    SB_LUT4 i1_3_lut_adj_173 (.I0(n4731), .I1(\lighthouse[0] ), .I2(n9989), 
            .I3(GND_net), .O(n23989));
    defparam i1_3_lut_adj_173.LUT_INIT = 16'h5454;
    SB_LUT4 Mux_34_i1_3_lut (.I0(ootx_payloads_0_241), .I1(ootx_payloads_1_241), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[241]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_34_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1808_5_lut (.I0(n2610), .I1(n2610), .I2(n2621), 
            .I3(n22679), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_17_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n22581), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_35_i1_3_lut (.I0(ootx_payloads_0_240), .I1(ootx_payloads_1_240), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[240]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_35_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1004_5 (.CI(n22457), .I0(n1410_c), .I1(n1433_c), 
            .CO(n22458));
    SB_CARRY mod_155_add_1473_17 (.CI(n22581), .I0(n2098), .I1(n2126), 
            .CO(n22582));
    SB_LUT4 i1_2_lut_adj_174 (.I0(\lighthouse[0] ), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n20098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i1_2_lut_adj_174.LUT_INIT = 16'h8888;
    SB_LUT4 Mux_36_i1_3_lut (.I0(ootx_payloads_0_239), .I1(ootx_payloads_1_239), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[239]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_36_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_175 (.I0(n109), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n1006));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_175.LUT_INIT = 16'h0080;
    SB_LUT4 i23_4_lut (.I0(n45_c), .I1(n3008), .I2(n40_adj_1908), .I3(n2989), 
            .O(n49_c));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n49_c), .I1(n47_c), .I2(n43_adj_1909), .I3(n44_c), 
            .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 Mux_21_i1_3_lut_adj_176 (.I0(data_counters_0_17), .I1(data_counters_1_17), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[17]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_21_i1_3_lut_adj_176.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_21_i1_3_lut_adj_177 (.I0(bit_counters_0_15), .I1(bit_counters_1_15), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[15]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_21_i1_3_lut_adj_177.LUT_INIT = 16'hcaca;
    SB_LUT4 i20509_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25177));
    defparam i20509_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 Mux_20_i1_3_lut_adj_178 (.I0(bit_counters_0_16), .I1(bit_counters_1_16), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[16]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_20_i1_3_lut_adj_178.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_179 (.I0(n109), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n750));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_179.LUT_INIT = 16'h0008;
    SB_LUT4 mod_155_add_1004_4_lut (.I0(n1411_c), .I1(n1411_c), .I2(n1433_c), 
            .I3(n22456), .O(n1510)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1808_5 (.CI(n22679), .I0(n2610), .I1(n2621), 
            .CO(n22680));
    SB_LUT4 mod_155_add_1473_16_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n22580), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1004_4 (.CI(n22456), .I0(n1411_c), .I1(n1433_c), 
            .CO(n22457));
    SB_LUT4 i7686_3_lut_4_lut (.I0(n888), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1250), .O(n11796));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7686_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_37_i1_3_lut (.I0(ootx_payloads_0_238), .I1(ootx_payloads_1_238), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[238]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_37_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1473_16 (.CI(n22580), .I0(n2099), .I1(n2126), 
            .CO(n22581));
    SB_LUT4 Mux_38_i1_3_lut (.I0(ootx_payloads_0_237), .I1(ootx_payloads_1_237), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[237]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_38_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1004_3_lut (.I0(n1412_c), .I1(n1412_c), .I2(n1433_c), 
            .I3(n22455), .O(n1511)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2076_24_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n22804), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2009_20_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n22772), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7094_3_lut_4_lut (.I0(n888), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_183), .O(n11204));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7094_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1942_13_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n22738), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_4_lut (.I0(n2611), .I1(n2611), .I2(n2621), 
            .I3(n22678), .O(n2710)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_15_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n22579), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1004_3 (.CI(n22455), .I0(n1412_c), .I1(n1433_c), 
            .CO(n22456));
    SB_LUT4 i1_2_lut_adj_180 (.I0(\lighthouse[0] ), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n112));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i1_2_lut_adj_180.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_181 (.I0(n119), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n888));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_181.LUT_INIT = 16'h0020;
    SB_CARRY mod_155_add_1473_15 (.CI(n22579), .I0(n2100), .I1(n2126), 
            .CO(n22580));
    SB_LUT4 mod_155_add_1004_2_lut (.I0(n2851[18]), .I1(n2851[18]), .I2(n25184), 
            .I3(VCC_net), .O(n1512)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1808_4 (.CI(n22678), .I0(n2611), .I1(n2621), 
            .CO(n22679));
    SB_LUT4 mod_155_add_1473_14_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n22578), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_182 (.I0(n119), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n632));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_182.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_1004_2 (.CI(VCC_net), .I0(n2851[18]), .I1(n25184), 
            .CO(n22455));
    SB_CARRY mod_155_add_1473_14 (.CI(n22578), .I0(n2101), .I1(n2126), 
            .CO(n22579));
    SB_LUT4 PrioSelect_105_i2_3_lut (.I0(data), .I1(n4485[5]), .I2(n34[1]), 
            .I3(GND_net), .O(n138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_105_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_937_14_lut (.I0(n1301_c), .I1(n1301_c), .I2(n1334_c), 
            .I3(n22454), .O(n1400_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1942_13 (.CI(n22738), .I0(n2802), .I1(n2819), 
            .CO(n22739));
    SB_LUT4 i7685_3_lut_4_lut (.I0(n886), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1251), .O(n11795));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7685_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1808_3_lut (.I0(n2612), .I1(n2612), .I2(n2621), 
            .I3(n22677), .O(n2711)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7093_3_lut_4_lut (.I0(n886), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_182), .O(n11203));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7093_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1473_13_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n22577), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_183 (.I0(n117), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n886));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_183.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_184 (.I0(n117), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n630));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_184.LUT_INIT = 16'h0002;
    SB_LUT4 i7549_3_lut_4_lut (.I0(n614), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1387), .O(n11659));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_937_13_lut (.I0(n1302_c), .I1(n1302_c), .I2(n1334_c), 
            .I3(n22453), .O(n1401_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_13 (.CI(n22577), .I0(n2102), .I1(n2126), 
            .CO(n22578));
    SB_LUT4 i1_4_lut_adj_185 (.I0(n3), .I1(n23993), .I2(n4729), .I3(n112), 
            .O(n23994));
    defparam i1_4_lut_adj_185.LUT_INIT = 16'hc8c0;
    SB_CARRY mod_155_add_937_13 (.CI(n22453), .I0(n1302_c), .I1(n1334_c), 
            .CO(n22454));
    SB_CARRY mod_155_add_1808_3 (.CI(n22677), .I0(n2612), .I1(n2621), 
            .CO(n22678));
    SB_LUT4 i1_3_lut_adj_186 (.I0(n22943), .I1(n23993), .I2(n4729), .I3(GND_net), 
            .O(n23996));
    defparam i1_3_lut_adj_186.LUT_INIT = 16'hc4c4;
    SB_LUT4 mod_155_add_1473_12_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n22576), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_937_12_lut (.I0(n1303_c), .I1(n1303_c), .I2(n1334_c), 
            .I3(n22452), .O(n1402_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7730_3_lut_4_lut (.I0(n976), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1206), .O(n11840));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7730_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_39_i1_3_lut (.I0(ootx_payloads_0_236), .I1(ootx_payloads_1_236), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[236]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_39_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7138_3_lut_4_lut (.I0(n976), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_227), .O(n11248));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7138_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1473_12 (.CI(n22576), .I0(n2103), .I1(n2126), 
            .CO(n22577));
    SB_CARRY mod_155_add_937_12 (.CI(n22452), .I0(n1303_c), .I1(n1334_c), 
            .CO(n22453));
    SB_LUT4 i6957_3_lut_4_lut (.I0(n614), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_46), .O(n11067));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6957_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2009_20 (.CI(n22772), .I0(n2895), .I1(n2918), 
            .CO(n22773));
    SB_LUT4 mod_155_add_1942_12_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n22737), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7684_3_lut_4_lut (.I0(n884), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1252), .O(n11794));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7684_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2143_32_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n22841), .O(n61_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_32_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1808_2_lut (.I0(n2851[6]), .I1(n2851[6]), .I2(n25178), 
            .I3(VCC_net), .O(n2712)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1473_11_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n22575), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_937_11_lut (.I0(n1304_c), .I1(n1304_c), .I2(n1334_c), 
            .I3(n22451), .O(n1403_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_11 (.CI(n22575), .I0(n2104), .I1(n2126), 
            .CO(n22576));
    SB_CARRY mod_155_add_2076_24 (.CI(n22804), .I0(n2991), .I1(n3017), 
            .CO(n22805));
    SB_CARRY mod_155_add_937_11 (.CI(n22451), .I0(n1304_c), .I1(n1334_c), 
            .CO(n22452));
    SB_CARRY mod_155_add_1808_2 (.CI(VCC_net), .I0(n2851[6]), .I1(n25178), 
            .CO(n22677));
    SB_LUT4 mod_155_add_1473_10_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n22574), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_937_10_lut (.I0(n1305_c), .I1(n1305_c), .I2(n1334_c), 
            .I3(n22450), .O(n1404_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_10 (.CI(n22574), .I0(n2105), .I1(n2126), 
            .CO(n22575));
    SB_LUT4 i7092_3_lut_4_lut (.I0(n884), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_181), .O(n11202));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7092_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_187 (.I0(n115), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n884));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_187.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_188 (.I0(n115), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n628));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_188.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_937_10 (.CI(n22450), .I0(n1305_c), .I1(n1334_c), 
            .CO(n22451));
    SB_LUT4 Mux_40_i1_3_lut (.I0(ootx_payloads_0_235), .I1(ootx_payloads_1_235), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[235]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_40_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1942_12 (.CI(n22737), .I0(n2803), .I1(n2819), 
            .CO(n22738));
    SB_LUT4 mod_155_add_1741_26_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n22676), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7683_3_lut_4_lut (.I0(n882), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1253), .O(n11793));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7683_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7091_3_lut_4_lut (.I0(n882), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_180), .O(n11201));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7091_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1473_9_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n22573), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_937_9_lut (.I0(n1306_c), .I1(n1306_c), .I2(n1334_c), 
            .I3(n22449), .O(n1405_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_41_i1_3_lut (.I0(ootx_payloads_0_234), .I1(ootx_payloads_1_234), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[234]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_41_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1473_9 (.CI(n22573), .I0(n2106), .I1(n2126), 
            .CO(n22574));
    SB_CARRY mod_155_add_937_9 (.CI(n22449), .I0(n1306_c), .I1(n1334_c), 
            .CO(n22450));
    SB_LUT4 mod_155_add_1741_25_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n22675), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_8_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n22572), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i110_2_lut_3_lut (.I0(n30_adj_1855), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n110_adj_1911));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i110_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mod_155_add_937_8_lut (.I0(n1307_c), .I1(n1307_c), .I2(n1334_c), 
            .I3(n22448), .O(n1406_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_8 (.CI(n22572), .I0(n2107), .I1(n2126), 
            .CO(n22573));
    SB_CARRY mod_155_add_937_8 (.CI(n22448), .I0(n1307_c), .I1(n1334_c), 
            .CO(n22449));
    SB_LUT4 i7578_3_lut_4_lut (.I0(n672), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1358), .O(n11688));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7578_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i109_2_lut_3_lut (.I0(n30_adj_1855), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i109_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY mod_155_add_2143_32 (.CI(n22841), .I0(n3084), .I1(n3116), 
            .CO(n22842));
    SB_LUT4 mod_155_add_2076_23_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n22803), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_3_lut_adj_189 (.I0(n4731), .I1(\lighthouse[0] ), .I2(n9989), 
            .I3(GND_net), .O(n23993));
    defparam i1_3_lut_adj_189.LUT_INIT = 16'h5151;
    SB_LUT4 i6986_3_lut_4_lut (.I0(n672), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_75), .O(n11096));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2009_19_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n22771), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_11_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n22736), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7548_3_lut_4_lut (.I0(n612), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1388), .O(n11658));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1741_25 (.CI(n22675), .I0(n2490), .I1(n2522), 
            .CO(n22676));
    SB_LUT4 mod_155_add_1473_7_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n22571), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6956_3_lut_4_lut (.I0(n612), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_45), .O(n11066));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6956_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_190 (.I0(n113), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n882));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_190.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_191 (.I0(n113), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n626));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_191.LUT_INIT = 16'h0002;
    SB_LUT4 i7682_3_lut_4_lut (.I0(n880), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1254), .O(n11792));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7682_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7090_3_lut_4_lut (.I0(n880), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_179), .O(n11200));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7090_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_192 (.I0(sensor_state_switch_counter[1]), .I1(sensor_state_switch_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_1914));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(32[9:36])
    defparam i1_2_lut_adj_192.LUT_INIT = 16'heeee;
    SB_LUT4 i7024_3_lut_4_lut (.I0(n748), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_113), .O(n11134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7024_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7616_3_lut_4_lut (.I0(n748), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1320), .O(n11726));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7616_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7729_3_lut_4_lut (.I0(n974), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1207), .O(n11839));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7729_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7137_3_lut_4_lut (.I0(n974), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_226), .O(n11247));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7137_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_193 (.I0(\lighthouse[0] ), .I1(n23993), .I2(n4729), 
            .I3(n23985), .O(n23995));
    defparam i1_4_lut_adj_193.LUT_INIT = 16'hc4c0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_194 (.I0(n111), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n880));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_194.LUT_INIT = 16'h0020;
    SB_LUT4 PrioSelect_101_i2_3_lut (.I0(data), .I1(n4485[4]), .I2(n34[1]), 
            .I3(GND_net), .O(n134));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_101_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_195 (.I0(n111), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n624));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_195.LUT_INIT = 16'h0002;
    SB_LUT4 PrioSelect_97_i2_3_lut (.I0(data), .I1(n4485[3]), .I2(n34[1]), 
            .I3(GND_net), .O(n130));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_97_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7681_3_lut_4_lut (.I0(n878), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1255), .O(n11791));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7681_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7089_3_lut_4_lut (.I0(n878), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_178), .O(n11199));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7089_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_196 (.I0(n107), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n1004));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_196.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_2143_31_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n22840), .O(n59_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_31_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_937_7_lut (.I0(n1308_c), .I1(n1308_c), .I2(n1334_c), 
            .I3(n22447), .O(n1407_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2009_19 (.CI(n22771), .I0(n2896), .I1(n2918), 
            .CO(n22772));
    SB_CARRY mod_155_add_1473_7 (.CI(n22571), .I0(n2108), .I1(n2126), 
            .CO(n22572));
    SB_CARRY mod_155_add_1942_11 (.CI(n22736), .I0(n2804), .I1(n2819), 
            .CO(n22737));
    SB_LUT4 PrioSelect_93_i2_3_lut (.I0(data), .I1(n4485[2]), .I2(n34[1]), 
            .I3(GND_net), .O(n126));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_93_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1741_24_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n22674), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut_adj_197 (.I0(sensor_state_switch_counter[4]), .I1(sensor_state_switch_counter[5]), 
            .I2(n37_adj_1914), .I3(sensor_state_switch_counter[3]), .O(n13329));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(32[9:36])
    defparam i1_4_lut_adj_197.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_198 (.I0(counter_from_last_rise_c[5]), .I1(counter_from_last_rise[4]), 
            .I2(GND_net), .I3(GND_net), .O(n291));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i1_2_lut_adj_198.LUT_INIT = 16'heeee;
    SB_LUT4 i19448_4_lut (.I0(\counter_from_last_rise[10] ), .I1(\counter_from_last_rise[9] ), 
            .I2(n22900), .I3(n4_adj_1917), .O(n24114));
    defparam i19448_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i19470_4_lut (.I0(\counter_from_last_rise[12] ), .I1(\counter_from_last_rise[11] ), 
            .I2(n9029), .I3(n24114), .O(data_N_1808));
    defparam i19470_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i11_4_lut_adj_199 (.I0(\counter_from_last_rise[21] ), .I1(\counter_from_last_rise[24] ), 
            .I2(\counter_from_last_rise[23] ), .I3(counter_from_last_rise[13]), 
            .O(n30_adj_1918));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(314[16:45])
    defparam i11_4_lut_adj_199.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_2076_23 (.CI(n22803), .I0(n2992), .I1(n3017), 
            .CO(n22804));
    SB_CARRY mod_155_add_937_7 (.CI(n22447), .I0(n1308_c), .I1(n1334_c), 
            .CO(n22448));
    SB_CARRY add_355_5 (.CI(n22277), .I0(counter_from_last_rise[3]), .I1(GND_net), 
            .CO(n22278));
    SB_LUT4 add_355_4_lut (.I0(GND_net), .I1(counter_from_last_rise[2]), 
            .I2(GND_net), .I3(n22276), .O(n6363)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1741_24 (.CI(n22674), .I0(n2491), .I1(n2522), 
            .CO(n22675));
    SB_LUT4 mod_155_add_1741_23_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n22673), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_4 (.CI(n22276), .I0(counter_from_last_rise[2]), .I1(GND_net), 
            .CO(n22277));
    SB_LUT4 mod_155_add_2009_18_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n22770), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_6_lut (.I0(n2109), .I1(n2109), .I2(n25185), 
            .I3(n22570), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_355_3_lut (.I0(GND_net), .I1(counter_from_last_rise[1]), 
            .I2(GND_net), .I3(n22275), .O(n6364)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1942_10_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n22735), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_937_6_lut (.I0(n1309_c), .I1(n1309_c), .I2(n25186), 
            .I3(n22446), .O(n1408_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1741_23 (.CI(n22673), .I0(n2492), .I1(n2522), 
            .CO(n22674));
    SB_CARRY add_355_3 (.CI(n22275), .I0(counter_from_last_rise[1]), .I1(GND_net), 
            .CO(n22276));
    SB_CARRY mod_155_add_1942_10 (.CI(n22735), .I0(n2805), .I1(n2819), 
            .CO(n22736));
    SB_CARRY mod_155_add_1473_6 (.CI(n22570), .I0(n2109), .I1(n25185), 
            .CO(n22571));
    SB_LUT4 add_154_4_lut (.I0(GND_net), .I1(n2849[2]), .I2(GND_net), 
            .I3(n22245), .O(n2851[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_154_4 (.CI(n22245), .I0(n2849[2]), .I1(GND_net), .CO(n22246));
    SB_CARRY mod_155_add_937_6 (.CI(n22446), .I0(n1309_c), .I1(n25186), 
            .CO(n22447));
    SB_LUT4 add_355_2_lut (.I0(GND_net), .I1(counter_from_last_rise[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n6365)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_154_3_lut (.I0(GND_net), .I1(n2849[1]), .I2(GND_net), 
            .I3(n22244), .O(n2851[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1741_22_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n22672), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_9_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n22734), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_12_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[10] ), 
            .I2(GND_net), .I3(n22223), .O(n337[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_66_12 (.CI(n22223), .I0(\ootx_payloads_N_1699[10] ), .I1(GND_net), 
            .CO(n22224));
    SB_CARRY mod_155_add_1741_22 (.CI(n22672), .I0(n2493), .I1(n2522), 
            .CO(n22673));
    SB_CARRY add_154_3 (.CI(n22244), .I0(n2849[1]), .I1(GND_net), .CO(n22245));
    SB_LUT4 mod_155_add_1741_21_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n22671), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1473_5_lut (.I0(n2110), .I1(n2110), .I2(n2126), 
            .I3(n22569), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_5 (.CI(n22569), .I0(n2110), .I1(n2126), 
            .CO(n22570));
    SB_CARRY add_355_2 (.CI(VCC_net), .I0(counter_from_last_rise[0]), .I1(GND_net), 
            .CO(n22275));
    SB_LUT4 add_154_2_lut (.I0(GND_net), .I1(n2849[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n2851[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_937_5_lut (.I0(n1310_c), .I1(n1310_c), .I2(n1334_c), 
            .I3(n22445), .O(n1409_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_2 (.CI(VCC_net), .I0(n2849[0]), .I1(GND_net), .CO(n22244));
    SB_LUT4 i15_4_lut_adj_200 (.I0(\counter_from_last_rise[26] ), .I1(n30_adj_1918), 
            .I2(\counter_from_last_rise[25] ), .I3(counter_from_last_rise[17]), 
            .O(n34_adj_1919));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(314[16:45])
    defparam i15_4_lut_adj_200.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_201 (.I0(\counter_from_last_rise[22] ), .I1(\counter_from_last_rise[31] ), 
            .I2(\counter_from_last_rise[29] ), .I3(counter_from_last_rise[14]), 
            .O(n32_adj_1920));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(314[16:45])
    defparam i13_4_lut_adj_201.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_202 (.I0(counter_from_last_rise[18]), .I1(\counter_from_last_rise[28] ), 
            .I2(\counter_from_last_rise[27] ), .I3(\counter_from_last_rise[30] ), 
            .O(n33_adj_1921));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(314[16:45])
    defparam i14_4_lut_adj_202.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_203 (.I0(counter_from_last_rise[15]), .I1(\counter_from_last_rise[19] ), 
            .I2(counter_from_last_rise[16]), .I3(\counter_from_last_rise[20] ), 
            .O(n31_adj_1922));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(314[16:45])
    defparam i12_4_lut_adj_203.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_204 (.I0(n31_adj_1922), .I1(n33_adj_1921), .I2(n32_adj_1920), 
            .I3(n34_adj_1919), .O(n9029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(314[16:45])
    defparam i18_4_lut_adj_204.LUT_INIT = 16'hfffe;
    SB_LUT4 i20311_4_lut (.I0(n24674), .I1(counter_from_last_rise[4]), .I2(\counter_from_last_rise[8] ), 
            .I3(counter_from_last_rise[3]), .O(n24679));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i20311_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i20310_4_lut (.I0(n24679), .I1(\counter_from_last_rise[6] ), 
            .I2(\counter_from_last_rise[8] ), .I3(counter_from_last_rise_c[5]), 
            .O(n24680));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i20310_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_205 (.I0(\counter_from_last_rise[9] ), .I1(n24680), 
            .I2(\counter_from_last_rise[8] ), .I3(\counter_from_last_rise[7] ), 
            .O(n271));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i1_4_lut_adj_205.LUT_INIT = 16'ha088;
    SB_LUT4 i15163_4_lut (.I0(\counter_from_last_rise[10] ), .I1(\counter_from_last_rise[12] ), 
            .I2(n271), .I3(\counter_from_last_rise[11] ), .O(n19257));
    defparam i15163_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 add_154_32_lut (.I0(GND_net), .I1(n2849[30]), .I2(GND_net), 
            .I3(n22273), .O(n2851[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_206 (.I0(n107), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n748));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_206.LUT_INIT = 16'h0008;
    SB_LUT4 mod_155_add_1473_4_lut (.I0(n2111), .I1(n2111), .I2(n2126), 
            .I3(n22568), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_4 (.CI(n22568), .I0(n2111), .I1(n2126), 
            .CO(n22569));
    SB_LUT4 add_66_32_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[30] ), 
            .I2(GND_net), .I3(n22243), .O(n337[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_66_11_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[9] ), 
            .I2(GND_net), .I3(n22222), .O(n337[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_937_5 (.CI(n22445), .I0(n1310_c), .I1(n1334_c), 
            .CO(n22446));
    SB_CARRY add_66_11 (.CI(n22222), .I0(\ootx_payloads_N_1699[9] ), .I1(GND_net), 
            .CO(n22223));
    SB_LUT4 add_66_31_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[29]), 
            .I2(GND_net), .I3(n22242), .O(n337[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_937_4_lut (.I0(n1311_adj_1923), .I1(n1311_adj_1923), 
            .I2(n1334_c), .I3(n22444), .O(n1410_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1741_21 (.CI(n22671), .I0(n2494), .I1(n2522), 
            .CO(n22672));
    SB_CARRY mod_155_add_2009_18 (.CI(n22770), .I0(n2897), .I1(n2918), 
            .CO(n22771));
    SB_CARRY mod_155_add_1942_9 (.CI(n22734), .I0(n2806), .I1(n2819), 
            .CO(n22735));
    SB_LUT4 mod_155_add_1473_3_lut (.I0(n2112), .I1(n2112), .I2(n2126), 
            .I3(n22567), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1741_20_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n22670), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_32 (.CI(n22273), .I0(n2849[30]), .I1(GND_net), .CO(n83));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_207 (.I0(n109), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n878));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_207.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_208 (.I0(n109), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n622));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_208.LUT_INIT = 16'h0002;
    SB_LUT4 Mux_42_i1_3_lut (.I0(ootx_payloads_0_233), .I1(ootx_payloads_1_233), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[233]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_42_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1741_20 (.CI(n22670), .I0(n2495), .I1(n2522), 
            .CO(n22671));
    SB_CARRY mod_155_add_937_4 (.CI(n22444), .I0(n1311_adj_1923), .I1(n1334_c), 
            .CO(n22445));
    SB_LUT4 add_154_31_lut (.I0(GND_net), .I1(n2849[29]), .I2(GND_net), 
            .I3(n22272), .O(n2851[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1741_19_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n22669), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1473_3 (.CI(n22567), .I0(n2112), .I1(n2126), 
            .CO(n22568));
    SB_CARRY add_154_31 (.CI(n22272), .I0(n2849[29]), .I1(GND_net), .CO(n22273));
    SB_LUT4 add_154_30_lut (.I0(GND_net), .I1(n2849[28]), .I2(GND_net), 
            .I3(n22271), .O(n2851[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1473_2_lut (.I0(n2851[11]), .I1(n2851[11]), .I2(n25185), 
            .I3(VCC_net), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_937_3_lut (.I0(n1312_adj_1925), .I1(n1312_adj_1925), 
            .I2(n1334_c), .I3(n22443), .O(n1411_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_8_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n22733), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1741_19 (.CI(n22669), .I0(n2496), .I1(n2522), 
            .CO(n22670));
    SB_LUT4 mod_155_add_2009_17_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n22769), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_30 (.CI(n22271), .I0(n2849[28]), .I1(GND_net), .CO(n22272));
    SB_CARRY add_66_31 (.CI(n22242), .I0(ootx_payloads_N_1699[29]), .I1(GND_net), 
            .CO(n22243));
    SB_CARRY mod_155_add_937_3 (.CI(n22443), .I0(n1312_adj_1925), .I1(n1334_c), 
            .CO(n22444));
    SB_LUT4 PrioSelect_89_i2_3_lut (.I0(data), .I1(n4485[1]), .I2(n34[1]), 
            .I3(GND_net), .O(n122));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_89_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1942_8 (.CI(n22733), .I0(n2807), .I1(n2819), 
            .CO(n22734));
    SB_LUT4 i1_2_lut_adj_209 (.I0(n13329), .I1(sensor_N_132), .I2(GND_net), 
            .I3(GND_net), .O(n6849));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(32[9:36])
    defparam i1_2_lut_adj_209.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_210 (.I0(sensor_state), .I1(data_N_1808), .I2(GND_net), 
            .I3(GND_net), .O(n23997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(199[5] 341[12])
    defparam i1_2_lut_adj_210.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_211 (.I0(counter_from_nskip_rise[18]), .I1(counter_from_nskip_rise[17]), 
            .I2(GND_net), .I3(GND_net), .O(n23967));
    defparam i1_2_lut_adj_211.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_212 (.I0(counter_from_nskip_rise[8]), .I1(counter_from_nskip_rise[6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1926));
    defparam i2_2_lut_adj_212.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_213 (.I0(counter_from_nskip_rise[4]), .I1(counter_from_nskip_rise[0]), 
            .I2(n7036), .I3(counter_from_nskip_rise[1]), .O(n22949));
    defparam i2_4_lut_adj_213.LUT_INIT = 16'hfefa;
    SB_LUT4 i3_4_lut_adj_214 (.I0(n22949), .I1(n6_adj_1926), .I2(counter_from_nskip_rise[7]), 
            .I3(counter_from_nskip_rise[5]), .O(n22878));
    defparam i3_4_lut_adj_214.LUT_INIT = 16'hfefc;
    SB_LUT4 i729_4_lut (.I0(counter_from_nskip_rise[10]), .I1(counter_from_nskip_rise[11]), 
            .I2(counter_from_nskip_rise[9]), .I3(n22878), .O(n24_adj_1927));
    defparam i729_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_4_lut_adj_215 (.I0(counter_from_nskip_rise[14]), .I1(counter_from_nskip_rise[13]), 
            .I2(n24_adj_1927), .I3(counter_from_nskip_rise[12]), .O(n22877));
    defparam i2_4_lut_adj_215.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_216 (.I0(n22877), .I1(n23967), .I2(counter_from_nskip_rise[16]), 
            .I3(counter_from_nskip_rise[15]), .O(n23970));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(260[9] 270[16])
    defparam i1_4_lut_adj_216.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_217 (.I0(n23997), .I1(n6849), .I2(n19257), .I3(n9029), 
            .O(n2280));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(199[5] 341[12])
    defparam i2_4_lut_adj_217.LUT_INIT = 16'h0008;
    SB_LUT4 add_66_30_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[28]), 
            .I2(GND_net), .I3(n22241), .O(n337[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_154_29_lut (.I0(GND_net), .I1(n2849[27]), .I2(GND_net), 
            .I3(n22270), .O(n2851[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1741_18_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n22668), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_30 (.CI(n22241), .I0(ootx_payloads_N_1699[28]), .I1(GND_net), 
            .CO(n22242));
    SB_LUT4 add_66_10_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[8] ), 
            .I2(GND_net), .I3(n22221), .O(n337[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1473_2 (.CI(VCC_net), .I0(n2851[11]), .I1(n25185), 
            .CO(n22567));
    SB_LUT4 mod_155_add_1406_21_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n22566), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_10 (.CI(n22221), .I0(\ootx_payloads_N_1699[8] ), .I1(GND_net), 
            .CO(n22222));
    SB_LUT4 add_66_29_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[27]), 
            .I2(GND_net), .I3(n22240), .O(n337[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_937_2_lut (.I0(n2851[19]), .I1(n2851[19]), .I2(n25186), 
            .I3(VCC_net), .O(n1412_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1741_18 (.CI(n22668), .I0(n2497), .I1(n2522), 
            .CO(n22669));
    SB_CARRY add_154_29 (.CI(n22270), .I0(n2849[27]), .I1(GND_net), .CO(n22271));
    SB_LUT4 i1_2_lut_adj_218 (.I0(\lighthouse[0] ), .I1(n4729), .I2(GND_net), 
            .I3(GND_net), .O(n23775));
    defparam i1_2_lut_adj_218.LUT_INIT = 16'h4444;
    SB_CARRY mod_155_add_937_2 (.CI(VCC_net), .I0(n2851[19]), .I1(n25186), 
            .CO(n22443));
    SB_LUT4 mod_155_add_1406_20_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n22565), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_29 (.CI(n22240), .I0(ootx_payloads_N_1699[27]), .I1(GND_net), 
            .CO(n22241));
    SB_LUT4 add_66_28_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[26]), 
            .I2(GND_net), .I3(n22239), .O(n337[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_870_13_lut (.I0(n1202_adj_1928), .I1(n1202_adj_1928), 
            .I2(n1235_c), .I3(n22442), .O(n1301_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_28_lut (.I0(GND_net), .I1(n2849[26]), .I2(GND_net), 
            .I3(n22269), .O(n2851[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_66_28 (.CI(n22239), .I0(ootx_payloads_N_1699[26]), .I1(GND_net), 
            .CO(n22240));
    SB_LUT4 mod_155_add_1942_7_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n22732), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1741_17_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n22667), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_9_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(GND_net), .I3(n22220), .O(n337[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_66_27_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[25]), 
            .I2(GND_net), .I3(n22238), .O(n337[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1406_20 (.CI(n22565), .I0(n1995), .I1(n2027), 
            .CO(n22566));
    SB_LUT4 mod_155_add_2076_22_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n22802), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2009_17 (.CI(n22769), .I0(n2898), .I1(n2918), 
            .CO(n22770));
    SB_CARRY mod_155_add_1741_17 (.CI(n22667), .I0(n2498), .I1(n2522), 
            .CO(n22668));
    SB_LUT4 mod_155_add_870_12_lut (.I0(n1203_adj_1929), .I1(n1203_adj_1929), 
            .I2(n1235_c), .I3(n22441), .O(n1302_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1942_7 (.CI(n22732), .I0(n2808), .I1(n2819), 
            .CO(n22733));
    SB_LUT4 mod_155_add_1741_16_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n22666), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1406_19_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n22564), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut_adj_219 (.I0(counter_from_nskip_rise[25]), .I1(counter_from_nskip_rise[27]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_1930));
    defparam i3_2_lut_adj_219.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_220 (.I0(counter_from_nskip_rise[28]), .I1(counter_from_nskip_rise[23]), 
            .I2(counter_from_nskip_rise[31]), .I3(counter_from_nskip_rise[24]), 
            .O(n22_adj_1931));
    defparam i9_4_lut_adj_220.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(counter_from_nskip_rise[22]), .I1(counter_from_nskip_rise[21]), 
            .I2(counter_from_nskip_rise[29]), .I3(GND_net), .O(n20_adj_1932));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_221 (.I0(counter_from_nskip_rise[19]), .I1(n22_adj_1931), 
            .I2(n16_adj_1930), .I3(counter_from_nskip_rise[20]), .O(n24_adj_1933));
    defparam i11_4_lut_adj_221.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_222 (.I0(counter_from_nskip_rise[26]), .I1(n24_adj_1933), 
            .I2(n20_adj_1932), .I3(counter_from_nskip_rise[30]), .O(n9196));
    defparam i12_4_lut_adj_222.LUT_INIT = 16'hfffe;
    SB_LUT4 i2961_2_lut (.I0(counter_from_nskip_rise[2]), .I1(counter_from_nskip_rise[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7036));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(260[13:45])
    defparam i2961_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_223 (.I0(counter_from_nskip_rise[6]), .I1(counter_from_nskip_rise[5]), 
            .I2(counter_from_nskip_rise[7]), .I3(n6_adj_1934), .O(n22857));
    defparam i4_4_lut_adj_223.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut_adj_224 (.I0(n22857), .I1(counter_from_nskip_rise[9]), 
            .I2(counter_from_nskip_rise[11]), .I3(counter_from_nskip_rise[10]), 
            .O(n10_adj_1935));
    defparam i4_4_lut_adj_224.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_225 (.I0(counter_from_nskip_rise[14]), .I1(counter_from_nskip_rise[16]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1936));
    defparam i2_2_lut_adj_225.LUT_INIT = 16'heeee;
    SB_CARRY add_154_28 (.CI(n22269), .I0(n2849[26]), .I1(GND_net), .CO(n22270));
    SB_LUT4 add_154_27_lut (.I0(GND_net), .I1(n2849[25]), .I2(GND_net), 
            .I3(n22268), .O(n2851[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1406_19 (.CI(n22564), .I0(n1996), .I1(n2027), 
            .CO(n22565));
    SB_CARRY mod_155_add_870_12 (.CI(n22441), .I0(n1203_adj_1929), .I1(n1235_c), 
            .CO(n22442));
    SB_CARRY mod_155_add_1741_16 (.CI(n22666), .I0(n2499), .I1(n2522), 
            .CO(n22667));
    SB_CARRY add_154_27 (.CI(n22268), .I0(n2849[25]), .I1(GND_net), .CO(n22269));
    SB_LUT4 mod_155_add_1942_6_lut (.I0(n2809), .I1(n2809), .I2(n25180), 
            .I3(n22731), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_154_26_lut (.I0(GND_net), .I1(n2849[24]), .I2(GND_net), 
            .I3(n22267), .O(n2851[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1942_6 (.CI(n22731), .I0(n2809), .I1(n25180), 
            .CO(n22732));
    SB_LUT4 i7680_3_lut_4_lut (.I0(n876), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1256), .O(n11790));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7680_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_870_11_lut (.I0(n1204_adj_1938), .I1(n1204_adj_1938), 
            .I2(n1235_c), .I3(n22440), .O(n1303_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1741_15_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n22665), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2143_31 (.CI(n22840), .I0(n3085), .I1(n3116), 
            .CO(n22841));
    SB_LUT4 mod_155_add_2143_30_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n22839), .O(n57_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_30_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1406_18_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n22563), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_43_i1_3_lut (.I0(ootx_payloads_0_232), .I1(ootx_payloads_1_232), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[232]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_43_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7088_3_lut_4_lut (.I0(n876), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_177), .O(n11198));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7088_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1406_18 (.CI(n22563), .I0(n1997), .I1(n2027), 
            .CO(n22564));
    SB_CARRY mod_155_add_870_11 (.CI(n22440), .I0(n1204_adj_1938), .I1(n1235_c), 
            .CO(n22441));
    SB_LUT4 i7547_3_lut_4_lut (.I0(n610), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1389), .O(n11657));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1406_17_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n22562), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2143_30 (.CI(n22839), .I0(n3086), .I1(n3116), 
            .CO(n22840));
    SB_LUT4 Mux_44_i1_3_lut (.I0(ootx_payloads_0_231), .I1(ootx_payloads_1_231), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[231]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_44_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_870_10_lut (.I0(n1205_adj_1940), .I1(n1205_adj_1940), 
            .I2(n1235_c), .I3(n22439), .O(n1304_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6955_3_lut_4_lut (.I0(n610), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_44), .O(n11065));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6955_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 PrioSelect_77_i2_3_lut (.I0(data), .I1(n4485[14]), .I2(n34[0]), 
            .I3(GND_net), .O(n110));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_77_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_226 (.I0(n107), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n876));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_226.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_227 (.I0(n107), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n620));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_227.LUT_INIT = 16'h0002;
    SB_LUT4 i7679_3_lut_4_lut (.I0(n874), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1257), .O(n11789));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7679_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7087_3_lut_4_lut (.I0(n874), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_176), .O(n11197));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7087_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7678_3_lut_4_lut (.I0(n872), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1258), .O(n11788));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7678_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7086_3_lut_4_lut (.I0(n872), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_175), .O(n11196));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7086_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i43_2_lut_3_lut (.I0(n20_adj_1943), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n43_adj_1944));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i43_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i76_2_lut_3_lut_4_lut (.I0(n20_adj_1943), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n76));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i76_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i75_2_lut_3_lut_4_lut (.I0(n20_adj_1943), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n75));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i75_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_228 (.I0(n103), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n872));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_228.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_229 (.I0(n103), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n616));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_229.LUT_INIT = 16'h0002;
    SB_LUT4 i7546_3_lut_4_lut (.I0(n608), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1390), .O(n11656));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6954_3_lut_4_lut (.I0(n608), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_43), .O(n11064));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6954_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7677_3_lut_4_lut (.I0(n870), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1259), .O(n11787));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7677_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7085_3_lut_4_lut (.I0(n870), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_174), .O(n11195));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7085_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7023_3_lut_4_lut (.I0(n746), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_112), .O(n11133));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7023_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7615_3_lut_4_lut (.I0(n746), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1321), .O(n11725));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7615_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7545_3_lut_4_lut (.I0(n606), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1391), .O(n11655));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6953_3_lut_4_lut (.I0(n606), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_42), .O(n11063));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6953_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_230 (.I0(n101), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n870));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_230.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_231 (.I0(n101), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n614));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_231.LUT_INIT = 16'h0002;
    SB_LUT4 i7544_3_lut_4_lut (.I0(n604), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1392), .O(n11654));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6952_3_lut_4_lut (.I0(n604), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_41), .O(n11062));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6952_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i234_2_lut_3_lut (.I0(n41_adj_1946), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n234));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i234_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i233_2_lut_3_lut (.I0(n41_adj_1946), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n233));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i233_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7005_3_lut_4_lut (.I0(n710), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_94), .O(n11115));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7597_3_lut_4_lut (.I0(n710), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1339), .O(n11707));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7597_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i41_2_lut_3_lut (.I0(n18_adj_1865), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n41_adj_1946));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i41_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i74_2_lut_3_lut_4_lut (.I0(n18_adj_1865), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n74_adj_1899));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i74_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i73_2_lut_3_lut_4_lut (.I0(n18_adj_1865), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n73));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i73_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_232 (.I0(n134_adj_1948), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n966));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_232.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_233 (.I0(n134_adj_1948), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n710));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_233.LUT_INIT = 16'h0008;
    SB_LUT4 i7676_3_lut_4_lut (.I0(n868), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1260), .O(n11786));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7676_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7084_3_lut_4_lut (.I0(n868), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_173), .O(n11194));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7084_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i134_2_lut_3_lut (.I0(n37_adj_1949), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n134_adj_1948));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i134_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i262_2_lut_3_lut_4_lut (.I0(n37_adj_1949), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n262));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i262_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 EnabledDecoder_2_i261_2_lut_3_lut_4_lut (.I0(n37_adj_1949), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n261));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i261_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7543_3_lut_4_lut (.I0(n602), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1393), .O(n11653));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6951_3_lut_4_lut (.I0(n602), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_40), .O(n11061));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6951_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_234 (.I0(n99), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n868));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_234.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_235 (.I0(n99), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n612));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_235.LUT_INIT = 16'h0002;
    SB_LUT4 i7022_3_lut_4_lut (.I0(n744), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_111), .O(n11132));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7022_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7614_3_lut_4_lut (.I0(n744), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1322), .O(n11724));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7614_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7675_3_lut_4_lut (.I0(n866), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1261), .O(n11785));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7675_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7083_3_lut_4_lut (.I0(n866), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_172), .O(n11193));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7083_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7542_3_lut_4_lut (.I0(n600), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1394), .O(n11652));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6885_3_lut_4_lut (.I0(n600), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_39), .O(n10995));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_236 (.I0(n103), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n1000));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_236.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_237 (.I0(n103), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n744));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_237.LUT_INIT = 16'h0008;
    SB_LUT4 i7674_3_lut_4_lut (.I0(n864), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1262), .O(n11784));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7674_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7082_3_lut_4_lut (.I0(n864), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_171), .O(n11192));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7082_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7541_3_lut_4_lut (.I0(n598), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1395), .O(n11651));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6910_3_lut_4_lut (.I0(n598), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_38), .O(n11020));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6910_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_45_i1_3_lut (.I0(ootx_payloads_0_230), .I1(ootx_payloads_1_230), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[230]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_45_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_46_i1_3_lut (.I0(ootx_payloads_0_229), .I1(ootx_payloads_1_229), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[229]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_46_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1741_15 (.CI(n22665), .I0(n2500), .I1(n2522), 
            .CO(n22666));
    SB_CARRY mod_155_add_870_10 (.CI(n22439), .I0(n1205_adj_1940), .I1(n1235_c), 
            .CO(n22440));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_238 (.I0(n95), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n864));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_238.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_239 (.I0(n95), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n608));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_239.LUT_INIT = 16'h0002;
    SB_LUT4 Mux_47_i1_3_lut (.I0(ootx_payloads_0_228), .I1(ootx_payloads_1_228), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[228]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_47_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_48_i1_3_lut (.I0(ootx_payloads_0_227), .I1(ootx_payloads_1_227), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[227]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_48_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7540_3_lut_4_lut (.I0(n596), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1396), .O(n11650));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7540_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6871_3_lut_4_lut (.I0(n596), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_37), .O(n10981));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6871_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7539_3_lut_4_lut (.I0(n594), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1397), .O(n11649));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7539_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_49_i1_3_lut (.I0(ootx_payloads_0_226), .I1(ootx_payloads_1_226), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[226]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_49_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_50_i1_3_lut (.I0(ootx_payloads_0_225), .I1(ootx_payloads_1_225), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[225]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_50_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1406_17 (.CI(n22562), .I0(n1998), .I1(n2027), 
            .CO(n22563));
    SB_LUT4 mod_155_add_1741_14_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n22664), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1741_14 (.CI(n22664), .I0(n2501), .I1(n2522), 
            .CO(n22665));
    SB_CARRY mod_155_add_2076_22 (.CI(n22802), .I0(n2993), .I1(n3017), 
            .CO(n22803));
    SB_LUT4 i6912_3_lut_4_lut (.I0(n594), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_36), .O(n11022));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6912_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_51_i1_3_lut (.I0(ootx_payloads_0_224), .I1(ootx_payloads_1_224), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[224]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_51_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i103_2_lut_3_lut (.I0(n39_adj_1902), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i103_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i168_2_lut_3_lut_4_lut (.I0(n39_adj_1902), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n168));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i168_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i252_2_lut_3_lut (.I0(n59_adj_1950), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n252));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i252_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i167_2_lut_3_lut_4_lut (.I0(n39_adj_1902), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n167));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i167_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i7538_3_lut_4_lut (.I0(n592), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1398), .O(n11648));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7538_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_adj_240 (.I0(n53_c), .I1(n13_adj_1951), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_1952));
    defparam i2_2_lut_adj_240.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_241 (.I0(n2851[0]), .I1(n3212), .I2(n3211), .I3(n3210), 
            .O(n22885));
    defparam i3_4_lut_adj_241.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_242 (.I0(n59_c), .I1(n25_adj_1953), .I2(n63_c), 
            .I3(n27_adj_1954), .O(n48_c));
    defparam i20_4_lut_adj_242.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_243 (.I0(n15_adj_1955), .I1(n33_adj_1956), .I2(n29_adj_1957), 
            .I3(n35_adj_1958), .O(n46_c));
    defparam i18_4_lut_adj_243.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_244 (.I0(n41_adj_1959), .I1(n47_adj_1960), .I2(n43_adj_1961), 
            .I3(n57_c), .O(n47_adj_1962));
    defparam i19_4_lut_adj_244.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_245 (.I0(n49_adj_1963), .I1(n61_c), .I2(n51_c), 
            .I3(n11), .O(n45_adj_1964));
    defparam i17_4_lut_adj_245.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_246 (.I0(n17_adj_1965), .I1(n37_adj_1966), .I2(n19_adj_1967), 
            .I3(n45_adj_1968), .O(n44_adj_1969));
    defparam i16_4_lut_adj_246.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_247 (.I0(n22885), .I1(n30_adj_1952), .I2(n21_adj_1970), 
            .I3(n3209), .O(n43_adj_1971));
    defparam i15_4_lut_adj_247.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45_adj_1964), .I1(n47_adj_1962), .I2(n46_c), 
            .I3(n48_c), .O(n54_c));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_248 (.I0(n31_adj_1972), .I1(n55_c), .I2(n39_adj_1973), 
            .I3(n23_adj_1974), .O(n49_adj_1975));
    defparam i21_4_lut_adj_248.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_1975), .I1(n54_c), .I2(n43_adj_1971), 
            .I3(n44_adj_1969), .O(n3215));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6870_3_lut_4_lut (.I0(n592), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_35), .O(n10980));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6870_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_52_i1_3_lut (.I0(ootx_payloads_0_223), .I1(ootx_payloads_1_223), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[223]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_52_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7021_3_lut_4_lut (.I0(n742), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_110), .O(n11131));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7021_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7613_3_lut_4_lut (.I0(n742), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1323), .O(n11723));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7613_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7673_3_lut_4_lut (.I0(n862), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1263), .O(n11783));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7673_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7081_3_lut_4_lut (.I0(n862), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_170), .O(n11191));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7081_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7537_3_lut_4_lut (.I0(n590), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1399), .O(n11647));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7537_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6875_3_lut_4_lut (.I0(n590), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_34), .O(n10985));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6875_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_53_i1_3_lut (.I0(ootx_payloads_0_222), .I1(ootx_payloads_1_222), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[222]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_53_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_54_i1_3_lut (.I0(ootx_payloads_0_221), .I1(ootx_payloads_1_221), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[221]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_54_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE i671__i2 (.Q(\ootx_payload_o[1][1] ), .C(clock_c), .E(n2283), 
            .D(n2[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_LUT4 Mux_55_i1_3_lut (.I0(ootx_payloads_0_220), .I1(ootx_payloads_1_220), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[220]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_55_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_56_i1_3_lut (.I0(ootx_payloads_0_219), .I1(ootx_payloads_1_219), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[219]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_56_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_57_i1_3_lut (.I0(ootx_payloads_0_218), .I1(ootx_payloads_1_218), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[218]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_57_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18191_3_lut (.I0(n3211), .I1(n3212), .I2(n2851[0]), .I3(GND_net), 
            .O(n6_adj_1977));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i18191_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i7536_3_lut_4_lut (.I0(n588), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1400), .O(n11646));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7536_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i18183_rep_10_2_lut (.I0(n3212), .I1(n2851[0]), .I2(GND_net), 
            .I3(GND_net), .O(n26307));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i18183_rep_10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_249 (.I0(n3211), .I1(n3210), .I2(n26307), .I3(n6_adj_1977), 
            .O(n6_adj_1979));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i2_4_lut_adj_249.LUT_INIT = 16'h1248;
    SB_LUT4 i18202_3_lut (.I0(n3209), .I1(n3210), .I2(n6_adj_1977), .I3(GND_net), 
            .O(n5328[4]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i18202_3_lut.LUT_INIT = 16'h5656;
    SB_LUT4 i19454_2_lut (.I0(n3209), .I1(n3212), .I2(GND_net), .I3(GND_net), 
            .O(n24120));
    defparam i19454_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20442_4_lut (.I0(n5328[4]), .I1(n6_adj_1979), .I2(n3212), 
            .I3(n2851[0]), .O(n24806));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i20442_4_lut.LUT_INIT = 16'h0440;
    SB_LUT4 i19477_4_lut (.I0(n3211), .I1(n3215), .I2(n3210), .I3(n24120), 
            .O(n24145));
    defparam i19477_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_250 (.I0(n24145), .I1(n24806), .I2(n2851[0]), 
            .I3(n3215), .O(n13));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[11:37])
    defparam i21_4_lut_adj_250.LUT_INIT = 16'hc505;
    SB_LUT4 Mux_58_i1_3_lut (.I0(ootx_payloads_0_217), .I1(ootx_payloads_1_217), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[217]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_58_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_870_9_lut (.I0(n1206_adj_1980), .I1(n1206_adj_1980), 
            .I2(n1235_c), .I3(n22438), .O(n1305_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1406_16_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n22561), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6890_3_lut_4_lut (.I0(n588), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_33), .O(n11000));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_59_i1_3_lut (.I0(ootx_payloads_0_216), .I1(ootx_payloads_1_216), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[216]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_59_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1406_16 (.CI(n22561), .I0(n1999), .I1(n2027), 
            .CO(n22562));
    SB_CARRY mod_155_add_870_9 (.CI(n22438), .I0(n1206_adj_1980), .I1(n1235_c), 
            .CO(n22439));
    SB_CARRY add_154_26 (.CI(n22267), .I0(n2849[24]), .I1(GND_net), .CO(n22268));
    SB_DFFE i671__i3 (.Q(\ootx_payload_o[1][2] ), .C(clock_c), .E(n2283), 
            .D(n2[2]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i4 (.Q(\ootx_payload_o[1][3] ), .C(clock_c), .E(n2283), 
            .D(n2[3]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i5 (.Q(\ootx_payload_o[1][4] ), .C(clock_c), .E(n2283), 
            .D(n2[4]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i6 (.Q(\ootx_payload_o[1][5] ), .C(clock_c), .E(n2283), 
            .D(n2[5]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i7 (.Q(\ootx_payload_o[1][6] ), .C(clock_c), .E(n2283), 
            .D(n2[6]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i8 (.Q(\ootx_payload_o[1][7] ), .C(clock_c), .E(n2283), 
            .D(n2[7]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i9 (.Q(\ootx_payload_o[1][8] ), .C(clock_c), .E(n2283), 
            .D(n2[8]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i10 (.Q(\ootx_payload_o[1][9] ), .C(clock_c), .E(n2283), 
            .D(n2[9]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i11 (.Q(\ootx_payload_o[1][10] ), .C(clock_c), .E(n2283), 
            .D(n2[10]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i12 (.Q(\ootx_payload_o[1][11] ), .C(clock_c), .E(n2283), 
            .D(n2[11]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i13 (.Q(\ootx_payload_o[1][12] ), .C(clock_c), .E(n2283), 
            .D(n2[12]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i14 (.Q(\ootx_payload_o[1][13] ), .C(clock_c), .E(n2283), 
            .D(n2[13]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i15 (.Q(\ootx_payload_o[1][14] ), .C(clock_c), .E(n2283), 
            .D(n2[14]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i16 (.Q(\ootx_payload_o[1][15] ), .C(clock_c), .E(n2283), 
            .D(n2[15]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i17 (.Q(\ootx_payload_o[1][16] ), .C(clock_c), .E(n2283), 
            .D(n2[16]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i18 (.Q(\ootx_payload_o[1][17] ), .C(clock_c), .E(n2283), 
            .D(n2[17]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i19 (.Q(\ootx_payload_o[1][18] ), .C(clock_c), .E(n2283), 
            .D(n2[18]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i20 (.Q(\ootx_payload_o[1][19] ), .C(clock_c), .E(n2283), 
            .D(n2[19]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i21 (.Q(\ootx_payload_o[1][20] ), .C(clock_c), .E(n2283), 
            .D(n2[20]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i22 (.Q(\ootx_payload_o[1][21] ), .C(clock_c), .E(n2283), 
            .D(n2[21]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i23 (.Q(\ootx_payload_o[1][22] ), .C(clock_c), .E(n2283), 
            .D(n2[22]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i24 (.Q(\ootx_payload_o[1][23] ), .C(clock_c), .E(n2283), 
            .D(n2[23]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i25 (.Q(\ootx_payload_o[1][24] ), .C(clock_c), .E(n2283), 
            .D(n2[24]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i26 (.Q(\ootx_payload_o[1][25] ), .C(clock_c), .E(n2283), 
            .D(n2[25]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i27 (.Q(\ootx_payload_o[1][26] ), .C(clock_c), .E(n2283), 
            .D(n2[26]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i28 (.Q(\ootx_payload_o[1][27] ), .C(clock_c), .E(n2283), 
            .D(n2[27]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i29 (.Q(\ootx_payload_o[1][28] ), .C(clock_c), .E(n2283), 
            .D(n2[28]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i30 (.Q(\ootx_payload_o[1][29] ), .C(clock_c), .E(n2283), 
            .D(n2[29]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i31 (.Q(\ootx_payload_o[1][30] ), .C(clock_c), .E(n2283), 
            .D(n2[30]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i32 (.Q(\ootx_payload_o[1][31] ), .C(clock_c), .E(n2283), 
            .D(n2[31]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i33 (.Q(\ootx_payload_o[1][32] ), .C(clock_c), .E(n2283), 
            .D(n2[32]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i34 (.Q(\ootx_payload_o[1][33] ), .C(clock_c), .E(n2283), 
            .D(n2[33]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i35 (.Q(\ootx_payload_o[1][34] ), .C(clock_c), .E(n2283), 
            .D(n2[34]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i36 (.Q(\ootx_payload_o[1][35] ), .C(clock_c), .E(n2283), 
            .D(n2[35]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i37 (.Q(\ootx_payload_o[1][36] ), .C(clock_c), .E(n2283), 
            .D(n2[36]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i38 (.Q(\ootx_payload_o[1][37] ), .C(clock_c), .E(n2283), 
            .D(n2[37]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i39 (.Q(\ootx_payload_o[1][38] ), .C(clock_c), .E(n2283), 
            .D(n2[38]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i40 (.Q(\ootx_payload_o[1][39] ), .C(clock_c), .E(n2283), 
            .D(n2[39]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i41 (.Q(\ootx_payload_o[1][40] ), .C(clock_c), .E(n2283), 
            .D(n2[40]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i42 (.Q(\ootx_payload_o[1][41] ), .C(clock_c), .E(n2283), 
            .D(n2[41]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i43 (.Q(\ootx_payload_o[1][42] ), .C(clock_c), .E(n2283), 
            .D(n2[42]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i44 (.Q(\ootx_payload_o[1][43] ), .C(clock_c), .E(n2283), 
            .D(n2[43]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i45 (.Q(\ootx_payload_o[1][44] ), .C(clock_c), .E(n2283), 
            .D(n2[44]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i46 (.Q(\ootx_payload_o[1][45] ), .C(clock_c), .E(n2283), 
            .D(n2[45]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i47 (.Q(\ootx_payload_o[1][46] ), .C(clock_c), .E(n2283), 
            .D(n2[46]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i48 (.Q(\ootx_payload_o[1][47] ), .C(clock_c), .E(n2283), 
            .D(n2[47]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i49 (.Q(\ootx_payload_o[1][48] ), .C(clock_c), .E(n2283), 
            .D(n2[48]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i50 (.Q(\ootx_payload_o[1][49] ), .C(clock_c), .E(n2283), 
            .D(n2[49]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i51 (.Q(\ootx_payload_o[1][50] ), .C(clock_c), .E(n2283), 
            .D(n2[50]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i52 (.Q(\ootx_payload_o[1][51] ), .C(clock_c), .E(n2283), 
            .D(n2[51]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i53 (.Q(\ootx_payload_o[1][52] ), .C(clock_c), .E(n2283), 
            .D(n2[52]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i54 (.Q(\ootx_payload_o[1][53] ), .C(clock_c), .E(n2283), 
            .D(n2[53]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i55 (.Q(\ootx_payload_o[1][54] ), .C(clock_c), .E(n2283), 
            .D(n2[54]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i56 (.Q(\ootx_payload_o[1][55] ), .C(clock_c), .E(n2283), 
            .D(n2[55]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i57 (.Q(\ootx_payload_o[1][56] ), .C(clock_c), .E(n2283), 
            .D(n2[56]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i58 (.Q(\ootx_payload_o[1][57] ), .C(clock_c), .E(n2283), 
            .D(n2[57]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i59 (.Q(\ootx_payload_o[1][58] ), .C(clock_c), .E(n2283), 
            .D(n2[58]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i60 (.Q(\ootx_payload_o[1][59] ), .C(clock_c), .E(n2283), 
            .D(n2[59]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i61 (.Q(\ootx_payload_o[1][60] ), .C(clock_c), .E(n2283), 
            .D(n2[60]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i62 (.Q(\ootx_payload_o[1][61] ), .C(clock_c), .E(n2283), 
            .D(n2[61]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i63 (.Q(\ootx_payload_o[1][62] ), .C(clock_c), .E(n2283), 
            .D(n2[62]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i64 (.Q(\ootx_payload_o[1][63] ), .C(clock_c), .E(n2283), 
            .D(n2[63]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i65 (.Q(\ootx_payload_o[1][64] ), .C(clock_c), .E(n2283), 
            .D(n2[64]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i66 (.Q(\ootx_payload_o[1][65] ), .C(clock_c), .E(n2283), 
            .D(n2[65]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i67 (.Q(\ootx_payload_o[1][66] ), .C(clock_c), .E(n2283), 
            .D(n2[66]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i68 (.Q(\ootx_payload_o[1][67] ), .C(clock_c), .E(n2283), 
            .D(n2[67]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i69 (.Q(\ootx_payload_o[1][68] ), .C(clock_c), .E(n2283), 
            .D(n2[68]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i70 (.Q(\ootx_payload_o[1][69] ), .C(clock_c), .E(n2283), 
            .D(n2[69]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i71 (.Q(\ootx_payload_o[1][70] ), .C(clock_c), .E(n2283), 
            .D(n2[70]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i72 (.Q(\ootx_payload_o[1][71] ), .C(clock_c), .E(n2283), 
            .D(n2[71]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i73 (.Q(\ootx_payload_o[1][72] ), .C(clock_c), .E(n2283), 
            .D(n2[72]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i74 (.Q(\ootx_payload_o[1][73] ), .C(clock_c), .E(n2283), 
            .D(n2[73]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i75 (.Q(\ootx_payload_o[1][74] ), .C(clock_c), .E(n2283), 
            .D(n2[74]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i76 (.Q(\ootx_payload_o[1][75] ), .C(clock_c), .E(n2283), 
            .D(n2[75]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i77 (.Q(\ootx_payload_o[1][76] ), .C(clock_c), .E(n2283), 
            .D(n2[76]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i78 (.Q(\ootx_payload_o[1][77] ), .C(clock_c), .E(n2283), 
            .D(n2[77]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i79 (.Q(\ootx_payload_o[1][78] ), .C(clock_c), .E(n2283), 
            .D(n2[78]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i80 (.Q(\ootx_payload_o[1][79] ), .C(clock_c), .E(n2283), 
            .D(n2[79]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i81 (.Q(\ootx_payload_o[1][80] ), .C(clock_c), .E(n2283), 
            .D(n2[80]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i82 (.Q(\ootx_payload_o[1][81] ), .C(clock_c), .E(n2283), 
            .D(n2[81]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i83 (.Q(\ootx_payload_o[1][82] ), .C(clock_c), .E(n2283), 
            .D(n2[82]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i84 (.Q(\ootx_payload_o[1][83] ), .C(clock_c), .E(n2283), 
            .D(n2[83]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i85 (.Q(\ootx_payload_o[1][84] ), .C(clock_c), .E(n2283), 
            .D(n2[84]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i86 (.Q(\ootx_payload_o[1][85] ), .C(clock_c), .E(n2283), 
            .D(n2[85]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i87 (.Q(\ootx_payload_o[1][86] ), .C(clock_c), .E(n2283), 
            .D(n2[86]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i88 (.Q(\ootx_payload_o[1][87] ), .C(clock_c), .E(n2283), 
            .D(n2[87]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i89 (.Q(\ootx_payload_o[1][88] ), .C(clock_c), .E(n2283), 
            .D(n2[88]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i90 (.Q(\ootx_payload_o[1][89] ), .C(clock_c), .E(n2283), 
            .D(n2[89]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i91 (.Q(\ootx_payload_o[1][90] ), .C(clock_c), .E(n2283), 
            .D(n2[90]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i92 (.Q(\ootx_payload_o[1][91] ), .C(clock_c), .E(n2283), 
            .D(n2[91]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i93 (.Q(\ootx_payload_o[1][92] ), .C(clock_c), .E(n2283), 
            .D(n2[92]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i94 (.Q(\ootx_payload_o[1][93] ), .C(clock_c), .E(n2283), 
            .D(n2[93]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i95 (.Q(\ootx_payload_o[1][94] ), .C(clock_c), .E(n2283), 
            .D(n2[94]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i96 (.Q(\ootx_payload_o[1][95] ), .C(clock_c), .E(n2283), 
            .D(n2[95]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i97 (.Q(\ootx_payload_o[1][96] ), .C(clock_c), .E(n2283), 
            .D(n2[96]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i98 (.Q(\ootx_payload_o[1][97] ), .C(clock_c), .E(n2283), 
            .D(n2[97]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i99 (.Q(\ootx_payload_o[1][98] ), .C(clock_c), .E(n2283), 
            .D(n2[98]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i100 (.Q(\ootx_payload_o[1][99] ), .C(clock_c), .E(n2283), 
            .D(n2[99]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i101 (.Q(\ootx_payload_o[1][100] ), .C(clock_c), .E(n2283), 
            .D(n2[100]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i102 (.Q(\ootx_payload_o[1][101] ), .C(clock_c), .E(n2283), 
            .D(n2[101]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i103 (.Q(\ootx_payload_o[1][102] ), .C(clock_c), .E(n2283), 
            .D(n2[102]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i104 (.Q(\ootx_payload_o[1][103] ), .C(clock_c), .E(n2283), 
            .D(n2[103]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i105 (.Q(\ootx_payload_o[1][104] ), .C(clock_c), .E(n2283), 
            .D(n2[104]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i106 (.Q(\ootx_payload_o[1][105] ), .C(clock_c), .E(n2283), 
            .D(n2[105]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i107 (.Q(\ootx_payload_o[1][106] ), .C(clock_c), .E(n2283), 
            .D(n2[106]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i108 (.Q(\ootx_payload_o[1][107] ), .C(clock_c), .E(n2283), 
            .D(n2[107]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i109 (.Q(\ootx_payload_o[1][108] ), .C(clock_c), .E(n2283), 
            .D(n2[108]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i110 (.Q(\ootx_payload_o[1][109] ), .C(clock_c), .E(n2283), 
            .D(n2[109]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i111 (.Q(\ootx_payload_o[1][110] ), .C(clock_c), .E(n2283), 
            .D(n2[110]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i112 (.Q(\ootx_payload_o[1][111] ), .C(clock_c), .E(n2283), 
            .D(n2[111]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i113 (.Q(\ootx_payload_o[1][112] ), .C(clock_c), .E(n2283), 
            .D(n2[112]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i114 (.Q(\ootx_payload_o[1][113] ), .C(clock_c), .E(n2283), 
            .D(n2[113]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i115 (.Q(\ootx_payload_o[1][114] ), .C(clock_c), .E(n2283), 
            .D(n2[114]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i116 (.Q(\ootx_payload_o[1][115] ), .C(clock_c), .E(n2283), 
            .D(n2[115]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i117 (.Q(\ootx_payload_o[1][116] ), .C(clock_c), .E(n2283), 
            .D(n2[116]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i118 (.Q(\ootx_payload_o[1][117] ), .C(clock_c), .E(n2283), 
            .D(n2[117]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i119 (.Q(\ootx_payload_o[1][118] ), .C(clock_c), .E(n2283), 
            .D(n2[118]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i120 (.Q(\ootx_payload_o[1][119] ), .C(clock_c), .E(n2283), 
            .D(n2[119]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i121 (.Q(\ootx_payload_o[1][120] ), .C(clock_c), .E(n2283), 
            .D(n2[120]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i122 (.Q(\ootx_payload_o[1][121] ), .C(clock_c), .E(n2283), 
            .D(n2[121]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i123 (.Q(\ootx_payload_o[1][122] ), .C(clock_c), .E(n2283), 
            .D(n2[122]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i124 (.Q(\ootx_payload_o[1][123] ), .C(clock_c), .E(n2283), 
            .D(n2[123]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i125 (.Q(\ootx_payload_o[1][124] ), .C(clock_c), .E(n2283), 
            .D(n2[124]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i126 (.Q(\ootx_payload_o[1][125] ), .C(clock_c), .E(n2283), 
            .D(n2[125]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i127 (.Q(\ootx_payload_o[1][126] ), .C(clock_c), .E(n2283), 
            .D(n2[126]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i128 (.Q(\ootx_payload_o[1][127] ), .C(clock_c), .E(n2283), 
            .D(n2[127]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i129 (.Q(\ootx_payload_o[1][128] ), .C(clock_c), .E(n2283), 
            .D(n2[128]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i130 (.Q(\ootx_payload_o[1][129] ), .C(clock_c), .E(n2283), 
            .D(n2[129]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i131 (.Q(\ootx_payload_o[1][130] ), .C(clock_c), .E(n2283), 
            .D(n2[130]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i132 (.Q(\ootx_payload_o[1][131] ), .C(clock_c), .E(n2283), 
            .D(n2[131]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i133 (.Q(\ootx_payload_o[1][132] ), .C(clock_c), .E(n2283), 
            .D(n2[132]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i134 (.Q(\ootx_payload_o[1][133] ), .C(clock_c), .E(n2283), 
            .D(n2[133]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i135 (.Q(\ootx_payload_o[1][134] ), .C(clock_c), .E(n2283), 
            .D(n2[134]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i136 (.Q(\ootx_payload_o[1][135] ), .C(clock_c), .E(n2283), 
            .D(n2[135]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i137 (.Q(\ootx_payload_o[1][136] ), .C(clock_c), .E(n2283), 
            .D(n2[136]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i138 (.Q(\ootx_payload_o[1][137] ), .C(clock_c), .E(n2283), 
            .D(n2[137]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i139 (.Q(\ootx_payload_o[1][138] ), .C(clock_c), .E(n2283), 
            .D(n2[138]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i140 (.Q(\ootx_payload_o[1][139] ), .C(clock_c), .E(n2283), 
            .D(n2[139]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i141 (.Q(\ootx_payload_o[1][140] ), .C(clock_c), .E(n2283), 
            .D(n2[140]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i142 (.Q(\ootx_payload_o[1][141] ), .C(clock_c), .E(n2283), 
            .D(n2[141]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i143 (.Q(\ootx_payload_o[1][142] ), .C(clock_c), .E(n2283), 
            .D(n2[142]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i144 (.Q(\ootx_payload_o[1][143] ), .C(clock_c), .E(n2283), 
            .D(n2[143]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i145 (.Q(\ootx_payload_o[1][144] ), .C(clock_c), .E(n2283), 
            .D(n2[144]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i146 (.Q(\ootx_payload_o[1][145] ), .C(clock_c), .E(n2283), 
            .D(n2[145]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i147 (.Q(\ootx_payload_o[1][146] ), .C(clock_c), .E(n2283), 
            .D(n2[146]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i148 (.Q(\ootx_payload_o[1][147] ), .C(clock_c), .E(n2283), 
            .D(n2[147]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i149 (.Q(\ootx_payload_o[1][148] ), .C(clock_c), .E(n2283), 
            .D(n2[148]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i150 (.Q(\ootx_payload_o[1][149] ), .C(clock_c), .E(n2283), 
            .D(n2[149]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i151 (.Q(\ootx_payload_o[1][150] ), .C(clock_c), .E(n2283), 
            .D(n2[150]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i152 (.Q(\ootx_payload_o[1][151] ), .C(clock_c), .E(n2283), 
            .D(n2[151]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i153 (.Q(\ootx_payload_o[1][152] ), .C(clock_c), .E(n2283), 
            .D(n2[152]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i154 (.Q(\ootx_payload_o[1][153] ), .C(clock_c), .E(n2283), 
            .D(n2[153]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i155 (.Q(\ootx_payload_o[1][154] ), .C(clock_c), .E(n2283), 
            .D(n2[154]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i156 (.Q(\ootx_payload_o[1][155] ), .C(clock_c), .E(n2283), 
            .D(n2[155]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i157 (.Q(\ootx_payload_o[1][156] ), .C(clock_c), .E(n2283), 
            .D(n2[156]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i158 (.Q(\ootx_payload_o[1][157] ), .C(clock_c), .E(n2283), 
            .D(n2[157]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i159 (.Q(\ootx_payload_o[1][158] ), .C(clock_c), .E(n2283), 
            .D(n2[158]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i160 (.Q(\ootx_payload_o[1][159] ), .C(clock_c), .E(n2283), 
            .D(n2[159]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i161 (.Q(\ootx_payload_o[1][160] ), .C(clock_c), .E(n2283), 
            .D(n2[160]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i162 (.Q(\ootx_payload_o[1][161] ), .C(clock_c), .E(n2283), 
            .D(n2[161]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i163 (.Q(\ootx_payload_o[1][162] ), .C(clock_c), .E(n2283), 
            .D(n2[162]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i164 (.Q(\ootx_payload_o[1][163] ), .C(clock_c), .E(n2283), 
            .D(n2[163]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i165 (.Q(\ootx_payload_o[1][164] ), .C(clock_c), .E(n2283), 
            .D(n2[164]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i166 (.Q(\ootx_payload_o[1][165] ), .C(clock_c), .E(n2283), 
            .D(n2[165]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i167 (.Q(\ootx_payload_o[1][166] ), .C(clock_c), .E(n2283), 
            .D(n2[166]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i168 (.Q(\ootx_payload_o[1][167] ), .C(clock_c), .E(n2283), 
            .D(n2[167]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i169 (.Q(\ootx_payload_o[1][168] ), .C(clock_c), .E(n2283), 
            .D(n2[168]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i170 (.Q(\ootx_payload_o[1][169] ), .C(clock_c), .E(n2283), 
            .D(n2[169]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i171 (.Q(\ootx_payload_o[1][170] ), .C(clock_c), .E(n2283), 
            .D(n2[170]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i172 (.Q(\ootx_payload_o[1][171] ), .C(clock_c), .E(n2283), 
            .D(n2[171]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i173 (.Q(\ootx_payload_o[1][172] ), .C(clock_c), .E(n2283), 
            .D(n2[172]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i174 (.Q(\ootx_payload_o[1][173] ), .C(clock_c), .E(n2283), 
            .D(n2[173]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i175 (.Q(\ootx_payload_o[1][174] ), .C(clock_c), .E(n2283), 
            .D(n2[174]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i176 (.Q(\ootx_payload_o[1][175] ), .C(clock_c), .E(n2283), 
            .D(n2[175]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i177 (.Q(\ootx_payload_o[1][176] ), .C(clock_c), .E(n2283), 
            .D(n2[176]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i178 (.Q(\ootx_payload_o[1][177] ), .C(clock_c), .E(n2283), 
            .D(n2[177]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i179 (.Q(\ootx_payload_o[1][178] ), .C(clock_c), .E(n2283), 
            .D(n2[178]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i180 (.Q(\ootx_payload_o[1][179] ), .C(clock_c), .E(n2283), 
            .D(n2[179]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i181 (.Q(\ootx_payload_o[1][180] ), .C(clock_c), .E(n2283), 
            .D(n2[180]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i182 (.Q(\ootx_payload_o[1][181] ), .C(clock_c), .E(n2283), 
            .D(n2[181]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i183 (.Q(\ootx_payload_o[1][182] ), .C(clock_c), .E(n2283), 
            .D(n2[182]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i184 (.Q(\ootx_payload_o[1][183] ), .C(clock_c), .E(n2283), 
            .D(n2[183]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i185 (.Q(\ootx_payload_o[1][184] ), .C(clock_c), .E(n2283), 
            .D(n2[184]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i186 (.Q(\ootx_payload_o[1][185] ), .C(clock_c), .E(n2283), 
            .D(n2[185]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i187 (.Q(\ootx_payload_o[1][186] ), .C(clock_c), .E(n2283), 
            .D(n2[186]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i188 (.Q(\ootx_payload_o[1][187] ), .C(clock_c), .E(n2283), 
            .D(n2[187]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i189 (.Q(\ootx_payload_o[1][188] ), .C(clock_c), .E(n2283), 
            .D(n2[188]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i190 (.Q(\ootx_payload_o[1][189] ), .C(clock_c), .E(n2283), 
            .D(n2[189]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i191 (.Q(\ootx_payload_o[1][190] ), .C(clock_c), .E(n2283), 
            .D(n2[190]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i192 (.Q(\ootx_payload_o[1][191] ), .C(clock_c), .E(n2283), 
            .D(n2[191]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i193 (.Q(\ootx_payload_o[1][192] ), .C(clock_c), .E(n2283), 
            .D(n2[192]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i194 (.Q(\ootx_payload_o[1][193] ), .C(clock_c), .E(n2283), 
            .D(n2[193]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i195 (.Q(\ootx_payload_o[1][194] ), .C(clock_c), .E(n2283), 
            .D(n2[194]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i196 (.Q(\ootx_payload_o[1][195] ), .C(clock_c), .E(n2283), 
            .D(n2[195]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i197 (.Q(\ootx_payload_o[1][196] ), .C(clock_c), .E(n2283), 
            .D(n2[196]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i198 (.Q(\ootx_payload_o[1][197] ), .C(clock_c), .E(n2283), 
            .D(n2[197]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i199 (.Q(\ootx_payload_o[1][198] ), .C(clock_c), .E(n2283), 
            .D(n2[198]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i200 (.Q(\ootx_payload_o[1][199] ), .C(clock_c), .E(n2283), 
            .D(n2[199]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i201 (.Q(\ootx_payload_o[1][200] ), .C(clock_c), .E(n2283), 
            .D(n2[200]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i202 (.Q(\ootx_payload_o[1][201] ), .C(clock_c), .E(n2283), 
            .D(n2[201]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i203 (.Q(\ootx_payload_o[1][202] ), .C(clock_c), .E(n2283), 
            .D(n2[202]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i204 (.Q(\ootx_payload_o[1][203] ), .C(clock_c), .E(n2283), 
            .D(n2[203]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i205 (.Q(\ootx_payload_o[1][204] ), .C(clock_c), .E(n2283), 
            .D(n2[204]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i206 (.Q(\ootx_payload_o[1][205] ), .C(clock_c), .E(n2283), 
            .D(n2[205]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i207 (.Q(\ootx_payload_o[1][206] ), .C(clock_c), .E(n2283), 
            .D(n2[206]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i208 (.Q(\ootx_payload_o[1][207] ), .C(clock_c), .E(n2283), 
            .D(n2[207]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i209 (.Q(\ootx_payload_o[1][208] ), .C(clock_c), .E(n2283), 
            .D(n2[208]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i210 (.Q(\ootx_payload_o[1][209] ), .C(clock_c), .E(n2283), 
            .D(n2[209]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i211 (.Q(\ootx_payload_o[1][210] ), .C(clock_c), .E(n2283), 
            .D(n2[210]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i212 (.Q(\ootx_payload_o[1][211] ), .C(clock_c), .E(n2283), 
            .D(n2[211]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i213 (.Q(\ootx_payload_o[1][212] ), .C(clock_c), .E(n2283), 
            .D(n2[212]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i214 (.Q(\ootx_payload_o[1][213] ), .C(clock_c), .E(n2283), 
            .D(n2[213]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i215 (.Q(\ootx_payload_o[1][214] ), .C(clock_c), .E(n2283), 
            .D(n2[214]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i216 (.Q(\ootx_payload_o[1][215] ), .C(clock_c), .E(n2283), 
            .D(n2[215]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i217 (.Q(\ootx_payload_o[1][216] ), .C(clock_c), .E(n2283), 
            .D(n2[216]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i218 (.Q(\ootx_payload_o[1][217] ), .C(clock_c), .E(n2283), 
            .D(n2[217]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i219 (.Q(\ootx_payload_o[1][218] ), .C(clock_c), .E(n2283), 
            .D(n2[218]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i220 (.Q(\ootx_payload_o[1][219] ), .C(clock_c), .E(n2283), 
            .D(n2[219]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i221 (.Q(\ootx_payload_o[1][220] ), .C(clock_c), .E(n2283), 
            .D(n2[220]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i222 (.Q(\ootx_payload_o[1][221] ), .C(clock_c), .E(n2283), 
            .D(n2[221]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i223 (.Q(\ootx_payload_o[1][222] ), .C(clock_c), .E(n2283), 
            .D(n2[222]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i224 (.Q(\ootx_payload_o[1][223] ), .C(clock_c), .E(n2283), 
            .D(n2[223]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i225 (.Q(\ootx_payload_o[1][224] ), .C(clock_c), .E(n2283), 
            .D(n2[224]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i226 (.Q(\ootx_payload_o[1][225] ), .C(clock_c), .E(n2283), 
            .D(n2[225]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i227 (.Q(\ootx_payload_o[1][226] ), .C(clock_c), .E(n2283), 
            .D(n2[226]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i228 (.Q(\ootx_payload_o[1][227] ), .C(clock_c), .E(n2283), 
            .D(n2[227]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i229 (.Q(\ootx_payload_o[1][228] ), .C(clock_c), .E(n2283), 
            .D(n2[228]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i230 (.Q(\ootx_payload_o[1][229] ), .C(clock_c), .E(n2283), 
            .D(n2[229]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i231 (.Q(\ootx_payload_o[1][230] ), .C(clock_c), .E(n2283), 
            .D(n2[230]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i232 (.Q(\ootx_payload_o[1][231] ), .C(clock_c), .E(n2283), 
            .D(n2[231]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i233 (.Q(\ootx_payload_o[1][232] ), .C(clock_c), .E(n2283), 
            .D(n2[232]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i234 (.Q(\ootx_payload_o[1][233] ), .C(clock_c), .E(n2283), 
            .D(n2[233]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i235 (.Q(\ootx_payload_o[1][234] ), .C(clock_c), .E(n2283), 
            .D(n2[234]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i236 (.Q(\ootx_payload_o[1][235] ), .C(clock_c), .E(n2283), 
            .D(n2[235]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i237 (.Q(\ootx_payload_o[1][236] ), .C(clock_c), .E(n2283), 
            .D(n2[236]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i238 (.Q(\ootx_payload_o[1][237] ), .C(clock_c), .E(n2283), 
            .D(n2[237]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i239 (.Q(\ootx_payload_o[1][238] ), .C(clock_c), .E(n2283), 
            .D(n2[238]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i240 (.Q(\ootx_payload_o[1][239] ), .C(clock_c), .E(n2283), 
            .D(n2[239]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i241 (.Q(\ootx_payload_o[1][240] ), .C(clock_c), .E(n2283), 
            .D(n2[240]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i242 (.Q(\ootx_payload_o[1][241] ), .C(clock_c), .E(n2283), 
            .D(n2[241]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i243 (.Q(\ootx_payload_o[1][242] ), .C(clock_c), .E(n2283), 
            .D(n2[242]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i244 (.Q(\ootx_payload_o[1][243] ), .C(clock_c), .E(n2283), 
            .D(n2[243]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i245 (.Q(\ootx_payload_o[1][244] ), .C(clock_c), .E(n2283), 
            .D(n2[244]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i246 (.Q(\ootx_payload_o[1][245] ), .C(clock_c), .E(n2283), 
            .D(n2[245]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i247 (.Q(\ootx_payload_o[1][246] ), .C(clock_c), .E(n2283), 
            .D(n2[246]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i248 (.Q(\ootx_payload_o[1][247] ), .C(clock_c), .E(n2283), 
            .D(n2[247]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i249 (.Q(\ootx_payload_o[1][248] ), .C(clock_c), .E(n2283), 
            .D(n2[248]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i250 (.Q(\ootx_payload_o[1][249] ), .C(clock_c), .E(n2283), 
            .D(n2[249]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i251 (.Q(\ootx_payload_o[1][250] ), .C(clock_c), .E(n2283), 
            .D(n2[250]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i252 (.Q(\ootx_payload_o[1][251] ), .C(clock_c), .E(n2283), 
            .D(n2[251]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i253 (.Q(\ootx_payload_o[1][252] ), .C(clock_c), .E(n2283), 
            .D(n2[252]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i254 (.Q(\ootx_payload_o[1][253] ), .C(clock_c), .E(n2283), 
            .D(n2[253]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i255 (.Q(\ootx_payload_o[1][254] ), .C(clock_c), .E(n2283), 
            .D(n2[254]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i256 (.Q(\ootx_payload_o[1][255] ), .C(clock_c), .E(n2283), 
            .D(n2[255]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i257 (.Q(\ootx_payload_o[1][256] ), .C(clock_c), .E(n2283), 
            .D(n2[256]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i258 (.Q(\ootx_payload_o[1][257] ), .C(clock_c), .E(n2283), 
            .D(n2[257]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i259 (.Q(\ootx_payload_o[1][258] ), .C(clock_c), .E(n2283), 
            .D(n2[258]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i260 (.Q(\ootx_payload_o[1][259] ), .C(clock_c), .E(n2283), 
            .D(n2[259]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i261 (.Q(\ootx_payload_o[1][260] ), .C(clock_c), .E(n2283), 
            .D(n2[260]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i262 (.Q(\ootx_payload_o[1][261] ), .C(clock_c), .E(n2283), 
            .D(n2[261]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i263 (.Q(\ootx_payload_o[1][262] ), .C(clock_c), .E(n2283), 
            .D(n2[262]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_DFFE i671__i264 (.Q(\ootx_payload_o[1][263] ), .C(clock_c), .E(n2283), 
            .D(n2[263]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_251 (.I0(n93_adj_2014), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n862));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_251.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_252 (.I0(n93_adj_2014), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n606));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_252.LUT_INIT = 16'h0002;
    SB_LUT4 i7672_3_lut_4_lut (.I0(n860), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1264), .O(n11782));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7672_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i932_933 (.Q(n1215), .C(clock_c), .D(n11831));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1406_15_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n22560), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2143_29_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n22838), .O(n55_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_5_lut (.I0(n2810), .I1(n2810), .I2(n2819), 
            .I3(n22730), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_870_8_lut (.I0(n1207_adj_2015), .I1(n1207_adj_2015), 
            .I2(n1235_c), .I3(n22437), .O(n1306_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2009_16_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n22768), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 PrioSelect_73_i2_3_lut (.I0(data), .I1(n4485[13]), .I2(n34[0]), 
            .I3(GND_net), .O(n106));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_73_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_60_i1_3_lut (.I0(ootx_payloads_0_215), .I1(ootx_payloads_1_215), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[215]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_60_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7080_3_lut_4_lut (.I0(n860), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_169), .O(n11190));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7080_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2009_16 (.CI(n22768), .I0(n2899), .I1(n2918), 
            .CO(n22769));
    SB_LUT4 i7535_3_lut_4_lut (.I0(n586), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1401), .O(n11645));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7535_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_61_i1_3_lut (.I0(ootx_payloads_0_214), .I1(ootx_payloads_1_214), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[214]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_61_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_870_8 (.CI(n22437), .I0(n1207_adj_2015), .I1(n1235_c), 
            .CO(n22438));
    SB_LUT4 mod_155_add_2076_21_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n22801), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2143_29 (.CI(n22838), .I0(n3087), .I1(n3116), 
            .CO(n22839));
    SB_LUT4 i6880_3_lut_4_lut (.I0(n586), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_32), .O(n10990));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6880_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2009_15_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n22767), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i251_2_lut_3_lut (.I0(n59_adj_1950), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n251));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i251_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_253 (.I0(n101), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n998));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_253.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_254 (.I0(n101), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n742));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_254.LUT_INIT = 16'h0008;
    SB_LUT4 i7577_3_lut_4_lut (.I0(n670), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1359), .O(n11687));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_62_i1_3_lut (.I0(ootx_payloads_0_213), .I1(ootx_payloads_1_213), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[213]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_62_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2009_15 (.CI(n22767), .I0(n2900), .I1(n2918), 
            .CO(n22768));
    SB_CARRY mod_155_add_1942_5 (.CI(n22730), .I0(n2810), .I1(n2819), 
            .CO(n22731));
    SB_LUT4 mod_155_add_1741_13_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n22663), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_4_lut (.I0(n2811), .I1(n2811), .I2(n2819), 
            .I3(n22729), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1406_15 (.CI(n22560), .I0(n2000), .I1(n2027), 
            .CO(n22561));
    SB_LUT4 mod_155_add_870_7_lut (.I0(n1208_adj_2017), .I1(n1208_adj_2017), 
            .I2(n1235_c), .I3(n22436), .O(n1307_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i101_2_lut_3_lut (.I0(n37_adj_1949), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i101_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 Mux_63_i1_3_lut (.I0(ootx_payloads_0_212), .I1(ootx_payloads_1_212), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[212]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_63_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i166_2_lut_3_lut_4_lut (.I0(n37_adj_1949), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n166_adj_2018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i166_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_1741_13 (.CI(n22663), .I0(n2502), .I1(n2522), 
            .CO(n22664));
    SB_LUT4 mod_155_add_1406_14_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n22559), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_38_i1_3_lut_adj_255 (.I0(data_counters_0_0), .I1(data_counters_1_0), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_38_i1_3_lut_adj_255.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_870_7 (.CI(n22436), .I0(n1208_adj_2017), .I1(n1235_c), 
            .CO(n22437));
    SB_LUT4 EnabledDecoder_2_i165_2_lut_3_lut_4_lut (.I0(n37_adj_1949), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n165));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i165_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 Mux_64_i1_3_lut (.I0(ootx_payloads_0_211), .I1(ootx_payloads_1_211), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[211]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_64_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 PrioSelect_69_i2_3_lut (.I0(data), .I1(n4485[12]), .I2(n34[0]), 
            .I3(GND_net), .O(n102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_69_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7534_3_lut_4_lut (.I0(n584), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1402), .O(n11644));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7534_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6985_3_lut_4_lut (.I0(n670), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_74), .O(n11095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6985_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1406_14 (.CI(n22559), .I0(n2001), .I1(n2027), 
            .CO(n22560));
    SB_LUT4 mod_155_add_1741_12_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n22662), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6907_3_lut_4_lut (.I0(n584), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_31), .O(n11017));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6907_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1406_13_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n22558), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7533_3_lut_4_lut (.I0(n582), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1403), .O(n11643));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7533_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6903_3_lut_4_lut (.I0(n582), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_30), .O(n11013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6903_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_65_i1_3_lut (.I0(ootx_payloads_0_210), .I1(ootx_payloads_1_210), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[210]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_65_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7671_3_lut_4_lut (.I0(n858), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1265), .O(n11781));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7671_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7079_3_lut_4_lut (.I0(n858), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_168), .O(n11189));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7079_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_66_i1_3_lut (.I0(ootx_payloads_0_209), .I1(ootx_payloads_1_209), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[209]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_66_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_870_6_lut (.I0(n1209_adj_2021), .I1(n1209_adj_2021), 
            .I2(n25189), .I3(n22435), .O(n1308_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_870_6 (.CI(n22435), .I0(n1209_adj_2021), .I1(n25189), 
            .CO(n22436));
    SB_LUT4 i7532_3_lut_4_lut (.I0(n580), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1404), .O(n11642));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 PrioSelect_65_i2_3_lut (.I0(data), .I1(n4485[11]), .I2(n34[0]), 
            .I3(GND_net), .O(n98));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_65_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1406_13 (.CI(n22558), .I0(n2002), .I1(n2027), 
            .CO(n22559));
    SB_LUT4 i6909_3_lut_4_lut (.I0(n580), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_29), .O(n11019));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6909_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1406_12_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n22557), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_870_5_lut (.I0(n1210_adj_2023), .I1(n1210_adj_2023), 
            .I2(n1235_c), .I3(n22434), .O(n1309_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1942_4 (.CI(n22729), .I0(n2811), .I1(n2819), 
            .CO(n22730));
    SB_LUT4 mod_155_add_2143_28_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n22837), .O(n53_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_67_i1_3_lut (.I0(ootx_payloads_0_208), .I1(ootx_payloads_1_208), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[208]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_67_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_870_5 (.CI(n22434), .I0(n1210_adj_2023), .I1(n1235_c), 
            .CO(n22435));
    SB_CARRY mod_155_add_1741_12 (.CI(n22662), .I0(n2503), .I1(n2522), 
            .CO(n22663));
    SB_LUT4 i7531_3_lut_4_lut (.I0(n578), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1405), .O(n11641));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2143_28 (.CI(n22837), .I0(n3088), .I1(n3116), 
            .CO(n22838));
    SB_LUT4 i7728_3_lut_4_lut (.I0(n972), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1208), .O(n11838));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7728_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6899_3_lut_4_lut (.I0(n578), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_28), .O(n11009));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6899_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1406_12 (.CI(n22557), .I0(n2003), .I1(n2027), 
            .CO(n22558));
    SB_LUT4 i7530_3_lut_4_lut (.I0(n576), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1406), .O(n11640));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7530_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_68_i1_3_lut (.I0(ootx_payloads_0_207), .I1(ootx_payloads_1_207), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[207]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_68_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_69_i1_3_lut (.I0(ootx_payloads_0_206), .I1(ootx_payloads_1_206), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[206]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_69_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6872_3_lut_4_lut (.I0(n576), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_27), .O(n10982));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6872_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_70_i1_3_lut (.I0(ootx_payloads_0_205), .I1(ootx_payloads_1_205), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[205]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_70_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_71_i1_3_lut (.I0(ootx_payloads_0_204), .I1(ootx_payloads_1_204), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[204]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_71_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2076_21 (.CI(n22801), .I0(n2994), .I1(n3017), 
            .CO(n22802));
    SB_LUT4 Mux_72_i1_3_lut (.I0(ootx_payloads_0_203), .I1(ootx_payloads_1_203), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[203]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_72_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7670_3_lut_4_lut (.I0(n856), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1266), .O(n11780));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7670_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7136_3_lut_4_lut (.I0(n972), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_225), .O(n11246));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7136_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2076_20_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n22800), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7078_3_lut_4_lut (.I0(n856), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_167), .O(n11188));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7078_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_73_i1_3_lut (.I0(ootx_payloads_0_202), .I1(ootx_payloads_1_202), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[202]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_73_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_2143_27_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n22836), .O(n51_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7529_3_lut_4_lut (.I0(n574), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1407), .O(n11639));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6873_3_lut_4_lut (.I0(n574), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_26), .O(n10983));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7727_3_lut_4_lut (.I0(n970), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1209), .O(n11837));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7727_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7135_3_lut_4_lut (.I0(n970), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_224), .O(n11245));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7135_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7726_3_lut_4_lut (.I0(n968), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1210), .O(n11836));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7726_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_256 (.I0(n87), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n856));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_256.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_257 (.I0(n87), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n600));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_257.LUT_INIT = 16'h0002;
    SB_LUT4 PrioSelect_61_i2_3_lut (.I0(data), .I1(n4485[10]), .I2(n34[0]), 
            .I3(GND_net), .O(n94));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_61_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7528_3_lut_4_lut (.I0(n572), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1408), .O(n11638));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7528_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6874_3_lut_4_lut (.I0(n572), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_25), .O(n10984));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6874_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_74_i1_3_lut (.I0(ootx_payloads_0_201), .I1(ootx_payloads_1_201), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[201]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_74_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7669_3_lut_4_lut (.I0(n854), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1267), .O(n11779));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7669_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7077_3_lut_4_lut (.I0(n854), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_166), .O(n11187));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7077_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15187_4_lut (.I0(counter_from_nskip_rise[8]), .I1(counter_from_nskip_rise[13]), 
            .I2(n10_adj_1935), .I3(counter_from_nskip_rise[12]), .O(n19283));
    defparam i15187_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 PrioSelect_57_i2_3_lut (.I0(data), .I1(n4485[9]), .I2(n34[0]), 
            .I3(GND_net), .O(n90));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_57_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7527_3_lut_4_lut (.I0(n570), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1409), .O(n11637));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7527_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7134_3_lut_4_lut (.I0(n968), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_223), .O(n11244));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7134_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6877_3_lut_4_lut (.I0(n570), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_24), .O(n10987));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6877_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7020_3_lut_4_lut (.I0(n740), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_109), .O(n11130));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7020_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7612_3_lut_4_lut (.I0(n740), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1324), .O(n11722));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7612_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_258 (.I0(n99), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n996));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_258.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_259 (.I0(n99), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n740));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_259.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i99_2_lut_3_lut (.I0(n35_adj_2030), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n99));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i99_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 Mux_75_i1_3_lut (.I0(ootx_payloads_0_200), .I1(ootx_payloads_1_200), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[200]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_75_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i164_2_lut_3_lut_4_lut (.I0(n35_adj_2030), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n164));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i164_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i163_2_lut_3_lut_4_lut (.I0(n35_adj_2030), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n163));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i163_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_260 (.I0(n85), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n854));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_260.LUT_INIT = 16'h0020;
    SB_LUT4 PrioSelect_53_i2_3_lut (.I0(data), .I1(n4485[8]), .I2(n34[0]), 
            .I3(GND_net), .O(n86));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_53_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_870_4_lut (.I0(n1211_adj_2031), .I1(n1211_adj_2031), 
            .I2(n1235_c), .I3(n22433), .O(n1310_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_261 (.I0(n85), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n598));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_261.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_2143_27 (.CI(n22836), .I0(n3089), .I1(n3116), 
            .CO(n22837));
    SB_LUT4 Mux_76_i1_3_lut (.I0(ootx_payloads_0_199), .I1(ootx_payloads_1_199), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[199]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_76_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7019_3_lut_4_lut (.I0(n738), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_108), .O(n11129));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7019_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1406_11_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n22556), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1741_11_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n22661), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 n25219_bdd_4_lut_4_lut (.I0(n35), .I1(ootx_payloads_N_1744[1]), 
            .I2(n13221), .I3(n25219), .O(n25222));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(94[10:59])
    defparam n25219_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i7611_3_lut_4_lut (.I0(n738), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1325), .O(n11721));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7611_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 PrioSelect_49_i2_3_lut (.I0(data), .I1(n4485[7]), .I2(n34[0]), 
            .I3(GND_net), .O(n82));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_49_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7526_3_lut_4_lut (.I0(n568), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1410), .O(n11636));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7526_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2143_26_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n22835), .O(n49_adj_1963)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_77_i1_3_lut (.I0(ootx_payloads_0_198), .I1(ootx_payloads_1_198), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[198]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_77_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6878_3_lut_4_lut (.I0(n568), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_23), .O(n10988));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7668_3_lut_4_lut (.I0(n852), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1268), .O(n11778));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7668_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_870_4 (.CI(n22433), .I0(n1211_adj_2031), .I1(n1235_c), 
            .CO(n22434));
    SB_LUT4 i7725_3_lut_4_lut (.I0(n966), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1211), .O(n11835));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7725_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2143_26 (.CI(n22835), .I0(n3090), .I1(n3116), 
            .CO(n22836));
    SB_CARRY mod_155_add_1741_11 (.CI(n22661), .I0(n2504), .I1(n2522), 
            .CO(n22662));
    SB_CARRY mod_155_add_1406_11 (.CI(n22556), .I0(n2004), .I1(n2027), 
            .CO(n22557));
    SB_CARRY mod_155_add_2076_20 (.CI(n22800), .I0(n2995), .I1(n3017), 
            .CO(n22801));
    SB_LUT4 i7076_3_lut_4_lut (.I0(n852), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_165), .O(n11186));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7076_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1406_10_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n22555), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i226_2_lut_3_lut (.I0(n66_adj_1904), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n226));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i226_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mod_155_add_870_3_lut (.I0(n1212_adj_2033), .I1(n1212_adj_2033), 
            .I2(n1235_c), .I3(n22432), .O(n1311_adj_1923)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_3_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_870_3 (.CI(n22432), .I0(n1212_adj_2033), .I1(n1235_c), 
            .CO(n22433));
    SB_LUT4 mod_155_add_2143_25_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n22834), .O(n47_adj_1960)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 PrioSelect_45_i2_3_lut (.I0(data), .I1(n4485[6]), .I2(n34[0]), 
            .I3(GND_net), .O(n78));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_45_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_78_i1_3_lut (.I0(ootx_payloads_0_197), .I1(ootx_payloads_1_197), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[197]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_78_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1406_10 (.CI(n22555), .I0(n2005), .I1(n2027), 
            .CO(n22556));
    SB_LUT4 mod_155_add_870_2_lut (.I0(n2851[20]), .I1(n2851[20]), .I2(n25189), 
            .I3(VCC_net), .O(n1312_adj_1925)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_4_lut_adj_262 (.I0(n19283), .I1(n23967), .I2(n6_adj_1936), 
            .I3(counter_from_nskip_rise[15]), .O(n23969));
    defparam i1_4_lut_adj_262.LUT_INIT = 16'hccc8;
    SB_LUT4 mod_155_add_1406_9_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n22554), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i225_2_lut_3_lut (.I0(n66_adj_1904), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n225));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i225_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY mod_155_add_870_2 (.CI(VCC_net), .I0(n2851[20]), .I1(n25189), 
            .CO(n22432));
    SB_LUT4 i7133_3_lut_4_lut (.I0(n966), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_222), .O(n11243));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7133_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7525_3_lut_4_lut (.I0(n566), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1411), .O(n11635));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1942_3_lut (.I0(n2812), .I1(n2812), .I2(n2819), 
            .I3(n22728), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1741_10_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n22660), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_79_i1_3_lut (.I0(ootx_payloads_0_196), .I1(ootx_payloads_1_196), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[196]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_79_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_80_i1_3_lut (.I0(ootx_payloads_0_195), .I1(ootx_payloads_1_195), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[195]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_80_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_81_i1_3_lut (.I0(ootx_payloads_0_194), .I1(ootx_payloads_1_194), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[194]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_81_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_66_27 (.CI(n22238), .I0(ootx_payloads_N_1699[25]), .I1(GND_net), 
            .CO(n22239));
    SB_LUT4 mod_155_add_2009_14_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n22766), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_26_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[24]), 
            .I2(GND_net), .I3(n22237), .O(n337[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_1406_9 (.CI(n22554), .I0(n2006), .I1(n2027), 
            .CO(n22555));
    SB_LUT4 i6879_3_lut_4_lut (.I0(n566), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_22), .O(n10989));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2076_19_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n22799), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_803_12_lut (.I0(n1103), .I1(n1103), .I2(n1136), 
            .I3(n22431), .O(n1202_adj_1928)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1942_3 (.CI(n22728), .I0(n2812), .I1(n2819), 
            .CO(n22729));
    SB_LUT4 Mux_82_i1_3_lut (.I0(ootx_payloads_0_193), .I1(ootx_payloads_1_193), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[193]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_82_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2076_19 (.CI(n22799), .I0(n2996), .I1(n3017), 
            .CO(n22800));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_263 (.I0(n83_adj_2035), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n852));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_263.LUT_INIT = 16'h0020;
    SB_CARRY mod_155_add_1741_10 (.CI(n22660), .I0(n2505), .I1(n2522), 
            .CO(n22661));
    SB_LUT4 mod_155_add_1942_2_lut (.I0(n2851[4]), .I1(n2851[4]), .I2(n25180), 
            .I3(VCC_net), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 Mux_83_i1_3_lut (.I0(ootx_payloads_0_192), .I1(ootx_payloads_1_192), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[192]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_83_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_264 (.I0(n83_adj_2035), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n596));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_264.LUT_INIT = 16'h0002;
    SB_LUT4 i7524_3_lut_4_lut (.I0(n564), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1412), .O(n11634));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2143_25 (.CI(n22834), .I0(n3091), .I1(n3116), 
            .CO(n22835));
    SB_LUT4 mod_155_add_2076_18_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n22798), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6881_3_lut_4_lut (.I0(n564), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_21), .O(n10991));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6881_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7667_3_lut_4_lut (.I0(n850), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1269), .O(n11777));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7667_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7075_3_lut_4_lut (.I0(n850), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_164), .O(n11185));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7075_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7576_3_lut_4_lut (.I0(n668), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1360), .O(n11686));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7523_3_lut_4_lut (.I0(n562), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1413), .O(n11633));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6882_3_lut_4_lut (.I0(n562), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_20), .O(n10992));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7004_3_lut_4_lut (.I0(n708), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_93), .O(n11114));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7004_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7596_3_lut_4_lut (.I0(n708), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1340), .O(n11706));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7596_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7522_3_lut_4_lut (.I0(n560), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1414), .O(n11632));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1406_8_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n22553), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1406_8 (.CI(n22553), .I0(n2007), .I1(n2027), 
            .CO(n22554));
    SB_LUT4 mod_155_add_803_11_lut (.I0(n1104), .I1(n1104), .I2(n1136), 
            .I3(n22430), .O(n1203_adj_1929)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_803_11 (.CI(n22430), .I0(n1104), .I1(n1136), 
            .CO(n22431));
    SB_LUT4 add_154_25_lut (.I0(GND_net), .I1(n2849[23]), .I2(GND_net), 
            .I3(n22266), .O(n2851[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6883_3_lut_4_lut (.I0(n560), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_19), .O(n10993));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6984_3_lut_4_lut (.I0(n668), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_73), .O(n11094));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6984_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_265 (.I0(n132), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n964));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_265.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_266 (.I0(n132), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n708));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_266.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_267 (.I0(n81), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n850));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_267.LUT_INIT = 16'h0020;
    SB_LUT4 mod_155_add_1741_9_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n22659), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1406_7_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n22552), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_26 (.CI(n22237), .I0(ootx_payloads_N_1699[24]), .I1(GND_net), 
            .CO(n22238));
    SB_CARRY mod_155_add_1741_9 (.CI(n22659), .I0(n2506), .I1(n2522), 
            .CO(n22660));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_268 (.I0(n81), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n594));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_268.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_1406_7 (.CI(n22552), .I0(n2008), .I1(n2027), 
            .CO(n22553));
    SB_LUT4 mod_155_add_803_10_lut (.I0(n1105), .I1(n1105), .I2(n1136), 
            .I3(n22429), .O(n1204_adj_1938)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_803_10 (.CI(n22429), .I0(n1105), .I1(n1136), 
            .CO(n22430));
    SB_LUT4 i3_4_lut_adj_269 (.I0(n9513), .I1(ootx_payloads_N_1698), .I2(n13), 
            .I3(n3), .O(ootx_payloads_N_1685));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i3_4_lut_adj_269.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i60_2_lut_3_lut (.I0(n20_adj_1943), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n60_adj_2038));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i60_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 Mux_37_i1_3_lut_adj_270 (.I0(data_counters_0_1), .I1(data_counters_1_1), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_37_i1_3_lut_adj_270.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i11_2_lut (.I0(ootx_payloads_N_1685), .I1(ootx_payloads_N_1699[0]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_2039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i11_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 Mux_36_i1_3_lut_adj_271 (.I0(data_counters_0_2), .I1(data_counters_1_2), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[2]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_36_i1_3_lut_adj_271.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i132_2_lut_3_lut (.I0(n35_adj_2030), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n132));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i132_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i260_2_lut_3_lut_4_lut (.I0(n35_adj_2030), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n260));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i260_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 EnabledDecoder_2_i259_2_lut_3_lut_4_lut (.I0(n35_adj_2030), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n259));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i259_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7521_3_lut_4_lut (.I0(n558), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1415), .O(n11631));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7521_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6884_3_lut_4_lut (.I0(n558), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_18), .O(n10994));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut (.I0(n20_adj_1943), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n59_adj_1950));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i59_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 PrioSelect_41_i2_3_lut (.I0(data), .I1(n4485[5]), .I2(n34[0]), 
            .I3(GND_net), .O(n74));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_41_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1741_8_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n22658), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_84_i1_3_lut (.I0(ootx_payloads_0_191), .I1(ootx_payloads_1_191), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[191]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_84_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1406_6_lut (.I0(n2009), .I1(n2009), .I2(n25188), 
            .I3(n22551), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1406_6 (.CI(n22551), .I0(n2009), .I1(n25188), 
            .CO(n22552));
    SB_CARRY add_66_9 (.CI(n22220), .I0(\ootx_payloads_N_1699[7] ), .I1(GND_net), 
            .CO(n22221));
    SB_LUT4 Mux_85_i1_3_lut (.I0(ootx_payloads_0_190), .I1(ootx_payloads_1_190), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[190]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_85_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_803_9_lut (.I0(n1106), .I1(n1106), .I2(n1136), 
            .I3(n22428), .O(n1205_adj_1940)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_803_9 (.CI(n22428), .I0(n1106), .I1(n1136), .CO(n22429));
    SB_LUT4 Mux_86_i1_3_lut (.I0(ootx_payloads_0_189), .I1(ootx_payloads_1_189), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[189]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_86_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_87_i1_3_lut (.I0(ootx_payloads_0_188), .I1(ootx_payloads_1_188), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[188]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_87_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_88_i1_3_lut (.I0(ootx_payloads_0_187), .I1(ootx_payloads_1_187), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[187]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_88_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2076_18 (.CI(n22798), .I0(n2997), .I1(n3017), 
            .CO(n22799));
    SB_LUT4 mod_155_add_1406_5_lut (.I0(n2010), .I1(n2010), .I2(n2027), 
            .I3(n22550), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2009_14 (.CI(n22766), .I0(n2901), .I1(n2918), 
            .CO(n22767));
    SB_CARRY mod_155_add_1942_2 (.CI(VCC_net), .I0(n2851[4]), .I1(n25180), 
            .CO(n22728));
    SB_LUT4 mod_155_add_803_8_lut (.I0(n1107), .I1(n1107), .I2(n1136), 
            .I3(n22427), .O(n1206_adj_1980)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_6_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(GND_net), .I3(n22217), .O(n337[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7666_3_lut_4_lut (.I0(n848), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1270), .O(n11776));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7666_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7074_3_lut_4_lut (.I0(n848), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_163), .O(n11184));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7074_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1741_8 (.CI(n22658), .I0(n2507), .I1(n2522), 
            .CO(n22659));
    SB_LUT4 mod_155_add_1875_28_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n22727), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_3_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[1]), .I2(GND_net), 
            .I3(n22214), .O(n337[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Mux_89_i1_3_lut (.I0(ootx_payloads_0_186), .I1(ootx_payloads_1_186), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[186]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_89_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7520_3_lut_4_lut (.I0(n556), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1416), .O(n11630));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7520_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1406_5 (.CI(n22550), .I0(n2010), .I1(n2027), 
            .CO(n22551));
    SB_LUT4 mod_155_add_1741_7_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n22657), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_90_i1_3_lut (.I0(ootx_payloads_0_185), .I1(ootx_payloads_1_185), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[185]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_90_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_91_i1_3_lut (.I0(ootx_payloads_0_184), .I1(ootx_payloads_1_184), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[184]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_91_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_803_8 (.CI(n22427), .I0(n1107), .I1(n1136), .CO(n22428));
    SB_LUT4 mod_155_add_1406_4_lut (.I0(n2011), .I1(n2011), .I2(n2027), 
            .I3(n22549), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_8_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(GND_net), .I3(n22219), .O(n337[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6886_3_lut_4_lut (.I0(n556), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_17), .O(n10996));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1406_4 (.CI(n22549), .I0(n2011), .I1(n2027), 
            .CO(n22550));
    SB_LUT4 mod_155_add_803_7_lut (.I0(n1108), .I1(n1108), .I2(n1136), 
            .I3(n22426), .O(n1207_adj_2015)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_25_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[23]), 
            .I2(GND_net), .I3(n22236), .O(n337[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_272 (.I0(n79), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n848));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_272.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_273 (.I0(n79), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n592));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_273.LUT_INIT = 16'h0002;
    SB_LUT4 Mux_35_i1_3_lut_adj_274 (.I0(data_counters_0_3), .I1(data_counters_1_3), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[3] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_35_i1_3_lut_adj_274.LUT_INIT = 16'hcaca;
    SB_LUT4 i7519_3_lut_4_lut (.I0(n554), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1417), .O(n11629));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6887_3_lut_4_lut (.I0(n554), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_16), .O(n10997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_803_7 (.CI(n22426), .I0(n1108), .I1(n1136), .CO(n22427));
    SB_LUT4 mod_155_add_1406_3_lut (.I0(n2012), .I1(n2012), .I2(n2027), 
            .I3(n22548), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 PrioSelect_37_i2_3_lut (.I0(data), .I1(n4485[4]), .I2(n34[0]), 
            .I3(GND_net), .O(n70));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_37_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1741_7 (.CI(n22657), .I0(n2508), .I1(n2522), 
            .CO(n22658));
    SB_LUT4 mod_155_add_803_6_lut (.I0(n1109), .I1(n1109), .I2(n25190), 
            .I3(n22425), .O(n1208_adj_2017)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1741_6_lut (.I0(n2509), .I1(n2509), .I2(n25187), 
            .I3(n22656), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 Mux_92_i1_3_lut (.I0(ootx_payloads_0_183), .I1(ootx_payloads_1_183), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[183]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_92_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7034_3_lut_4_lut (.I0(n768), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_123), .O(n11144));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7034_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1406_3 (.CI(n22548), .I0(n2012), .I1(n2027), 
            .CO(n22549));
    SB_LUT4 i7626_3_lut_4_lut (.I0(n768), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1310), .O(n11736));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7626_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7665_3_lut_4_lut (.I0(n846), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1271), .O(n11775));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7665_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_803_6 (.CI(n22425), .I0(n1109), .I1(n25190), 
            .CO(n22426));
    SB_CARRY mod_155_add_1741_6 (.CI(n22656), .I0(n2509), .I1(n25187), 
            .CO(n22657));
    SB_LUT4 Mux_93_i1_3_lut (.I0(ootx_payloads_0_182), .I1(ootx_payloads_1_182), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[182]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_93_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1406_2_lut (.I0(n2851[12]), .I1(n2851[12]), .I2(n25188), 
            .I3(VCC_net), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1406_2 (.CI(VCC_net), .I0(n2851[12]), .I1(n25188), 
            .CO(n22548));
    SB_CARRY add_154_25 (.CI(n22266), .I0(n2849[23]), .I1(GND_net), .CO(n22267));
    SB_LUT4 i7073_3_lut_4_lut (.I0(n846), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_162), .O(n11183));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7073_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_275 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n92), .O(n540));
    defparam i1_2_lut_3_lut_4_lut_adj_275.LUT_INIT = 16'h0100;
    SB_LUT4 mod_155_add_803_5_lut (.I0(n1110), .I1(n1110), .I2(n1136), 
            .I3(n22424), .O(n1209_adj_2021)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_803_5 (.CI(n22424), .I0(n1110), .I1(n1136), .CO(n22425));
    SB_CARRY add_66_25 (.CI(n22236), .I0(ootx_payloads_N_1699[23]), .I1(GND_net), 
            .CO(n22237));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_276 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n94_adj_1872), .O(n542));
    defparam i1_2_lut_3_lut_4_lut_adj_276.LUT_INIT = 16'h0100;
    SB_LUT4 mod_155_add_1875_27_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n22726), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1339_20_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n22547), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_24_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[22]), 
            .I2(GND_net), .I3(n22235), .O(n337[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_277 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n96), .O(n544));
    defparam i1_2_lut_3_lut_4_lut_adj_277.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_278 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n110_adj_1911), .O(n558));
    defparam i1_2_lut_3_lut_4_lut_adj_278.LUT_INIT = 16'h0100;
    SB_LUT4 mod_155_add_1741_5_lut (.I0(n2510), .I1(n2510), .I2(n2522), 
            .I3(n22655), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_803_4_lut (.I0(n1111), .I1(n1111), .I2(n1136), 
            .I3(n22423), .O(n1210_adj_2023)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_154_24_lut (.I0(GND_net), .I1(n2849[22]), .I2(GND_net), 
            .I3(n22265), .O(n2851[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_279 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n162_adj_1905), .I3(GND_net), .O(n546));
    defparam i1_2_lut_3_lut_adj_279.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_280 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n164), .I3(GND_net), .O(n548));
    defparam i1_2_lut_3_lut_adj_280.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1339_19_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n22546), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2143_24_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n22833), .O(n45_adj_1968)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut_4_lut (.I0(n11_adj_2039), .I1(ootx_payloads_N_1699[1]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(ootx_payloads_N_1699[2]), 
            .O(n35_adj_2030));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i35_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY mod_155_add_803_4 (.CI(n22423), .I0(n1111), .I1(n1136), .CO(n22424));
    SB_LUT4 mod_155_add_2076_17_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n22797), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_24 (.CI(n22235), .I0(ootx_payloads_N_1699[22]), .I1(GND_net), 
            .CO(n22236));
    SB_LUT4 Mux_94_i1_3_lut (.I0(ootx_payloads_0_181), .I1(ootx_payloads_1_181), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[181]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_94_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_281 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n166_adj_2018), .I3(GND_net), .O(n550));
    defparam i1_2_lut_3_lut_adj_281.LUT_INIT = 16'h1010;
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut_4_lut (.I0(n11_adj_2039), .I1(ootx_payloads_N_1699[1]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(ootx_payloads_N_1699[2]), 
            .O(n36_adj_2041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i36_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_CARRY mod_155_add_1339_19 (.CI(n22546), .I0(n1896), .I1(n1928), 
            .CO(n22547));
    SB_LUT4 mod_155_add_2009_13_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n22765), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_8 (.CI(n22219), .I0(\ootx_payloads_N_1699[6] ), .I1(GND_net), 
            .CO(n22220));
    SB_LUT4 i1_2_lut_3_lut_adj_282 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n168), .I3(GND_net), .O(n552));
    defparam i1_2_lut_3_lut_adj_282.LUT_INIT = 16'h1010;
    SB_LUT4 i7566_3_lut_4_lut (.I0(n648), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1370), .O(n11676));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_283 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n170_adj_2042), .I3(GND_net), .O(n554));
    defparam i1_2_lut_3_lut_adj_283.LUT_INIT = 16'h1010;
    SB_LUT4 i15158_4_lut (.I0(n9196), .I1(n2280), .I2(n23970), .I3(n23969), 
            .O(n19251));
    defparam i15158_4_lut.LUT_INIT = 16'hc8cc;
    SB_LUT4 mod_155_add_803_3_lut (.I0(n1112), .I1(n1112), .I2(n1136), 
            .I3(n22422), .O(n1211_adj_2031)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_3_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_27 (.CI(n22726), .I0(n2688), .I1(n2720), 
            .CO(n22727));
    SB_CARRY mod_155_add_1741_5 (.CI(n22655), .I0(n2510), .I1(n2522), 
            .CO(n22656));
    SB_LUT4 mod_155_add_1741_4_lut (.I0(n2511), .I1(n2511), .I2(n2522), 
            .I3(n22654), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_adj_284 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n172), .I3(GND_net), .O(n556));
    defparam i1_2_lut_3_lut_adj_284.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_285 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n112_adj_2043), .O(n560));
    defparam i1_2_lut_3_lut_4_lut_adj_285.LUT_INIT = 16'h0100;
    SB_LUT4 i6974_3_lut_4_lut (.I0(n648), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_63), .O(n11084));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6974_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1339_18_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n22545), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_18 (.CI(n22545), .I0(n1897), .I1(n1928), 
            .CO(n22546));
    SB_CARRY add_66_3 (.CI(n22214), .I0(ootx_payloads_N_1699[1]), .I1(GND_net), 
            .CO(n22215));
    SB_CARRY mod_155_add_803_3 (.CI(n22422), .I0(n1112), .I1(n1136), .CO(n22423));
    SB_LUT4 mod_155_add_803_2_lut (.I0(n2851[21]), .I1(n2851[21]), .I2(n25190), 
            .I3(VCC_net), .O(n1212_adj_2033)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_66_7_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(n22218), .O(n337[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_286 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n95), .O(n736));
    defparam i1_2_lut_3_lut_4_lut_adj_286.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_287 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n110_adj_1911), .O(n686));
    defparam i1_2_lut_3_lut_4_lut_adj_287.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_1339_17_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n22544), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_17 (.CI(n22544), .I0(n1898), .I1(n1928), 
            .CO(n22545));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_288 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n114_adj_2044), .O(n690));
    defparam i1_2_lut_3_lut_4_lut_adj_288.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_95_i1_3_lut (.I0(ootx_payloads_0_180), .I1(ootx_payloads_1_180), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[180]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_95_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_803_2 (.CI(VCC_net), .I0(n2851[21]), .I1(n25190), 
            .CO(n22422));
    SB_LUT4 i7031_3_lut_4_lut (.I0(n762), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_120), .O(n11141));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7031_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_289 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n116), .O(n692));
    defparam i1_2_lut_3_lut_4_lut_adj_289.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_96_i1_3_lut (.I0(ootx_payloads_0_179), .I1(ootx_payloads_1_179), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[179]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_96_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2009_13 (.CI(n22765), .I0(n2902), .I1(n2918), 
            .CO(n22766));
    SB_LUT4 mod_155_add_736_11_lut (.I0(n1004_c), .I1(n1004_c), .I2(n1037), 
            .I3(n22421), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_23_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[21]), 
            .I2(GND_net), .I3(n22234), .O(n337[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1875_26_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n22725), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1741_4 (.CI(n22654), .I0(n2511), .I1(n2522), 
            .CO(n22655));
    SB_LUT4 mod_155_add_2009_12_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n22764), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7623_3_lut_4_lut (.I0(n762), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1313), .O(n11733));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7623_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_290 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n120), .O(n696));
    defparam i1_2_lut_3_lut_4_lut_adj_290.LUT_INIT = 16'h1000;
    SB_LUT4 EnabledDecoder_2_i250_2_lut_3_lut (.I0(n57_adj_2045), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n250));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i250_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i249_2_lut_3_lut (.I0(n57_adj_2045), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n249));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i249_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_291 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n122_adj_2046), .O(n698));
    defparam i1_2_lut_3_lut_4_lut_adj_291.LUT_INIT = 16'h1000;
    SB_LUT4 lighthouse_counter_639_mux_6_i1_4_lut (.I0(n129[0]), .I1(n9196), 
            .I2(n19251), .I3(n23970), .O(n69[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam lighthouse_counter_639_mux_6_i1_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 mod_155_add_1741_3_lut (.I0(n2512), .I1(n2512), .I2(n2522), 
            .I3(n22653), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1339_16_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n22543), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_97_i1_3_lut (.I0(ootx_payloads_0_178), .I1(ootx_payloads_1_178), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[178]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_97_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_292 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n124), .O(n700));
    defparam i1_2_lut_3_lut_4_lut_adj_292.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_293 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n128), .O(n576));
    defparam i1_2_lut_3_lut_4_lut_adj_293.LUT_INIT = 16'h0100;
    SB_CARRY mod_155_add_1339_16 (.CI(n22543), .I0(n1899), .I1(n1928), 
            .CO(n22544));
    SB_LUT4 mod_155_add_736_10_lut (.I0(n1005), .I1(n1005), .I2(n1037), 
            .I3(n22420), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_26 (.CI(n22725), .I0(n2689), .I1(n2720), 
            .CO(n22726));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_294 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n126_adj_1853), .O(n702));
    defparam i1_2_lut_3_lut_4_lut_adj_294.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_98_i1_3_lut (.I0(ootx_payloads_0_177), .I1(ootx_payloads_1_177), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[177]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_98_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7710_3_lut_4_lut (.I0(n936), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1226), .O(n11820));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7710_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_99_i1_3_lut (.I0(ootx_payloads_0_176), .I1(ootx_payloads_1_176), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[176]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_99_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_736_10 (.CI(n22420), .I0(n1005), .I1(n1037), 
            .CO(n22421));
    SB_LUT4 mod_155_add_1339_15_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n22542), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1741_3 (.CI(n22653), .I0(n2512), .I1(n2522), 
            .CO(n22654));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_295 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n128), .O(n704));
    defparam i1_2_lut_3_lut_4_lut_adj_295.LUT_INIT = 16'h1000;
    SB_LUT4 i7724_3_lut_4_lut (.I0(n964), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1212), .O(n11834));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7724_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_296 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n136), .O(n584));
    defparam i1_2_lut_3_lut_4_lut_adj_296.LUT_INIT = 16'h0100;
    SB_LUT4 Mux_100_i1_3_lut (.I0(ootx_payloads_0_175), .I1(ootx_payloads_1_175), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[175]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_100_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1339_15 (.CI(n22542), .I0(n1900), .I1(n1928), 
            .CO(n22543));
    SB_LUT4 mod_155_add_736_9_lut (.I0(n1006_c), .I1(n1006_c), .I2(n1037), 
            .I3(n22419), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_736_9 (.CI(n22419), .I0(n1006_c), .I1(n1037), 
            .CO(n22420));
    SB_LUT4 Mux_101_i1_3_lut (.I0(ootx_payloads_0_174), .I1(ootx_payloads_1_174), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[174]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_101_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_297 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n130_adj_2047), .O(n706));
    defparam i1_2_lut_3_lut_4_lut_adj_297.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_1741_2_lut (.I0(n2851[7]), .I1(n2851[7]), .I2(n25187), 
            .I3(VCC_net), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1875_25_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n22724), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_24 (.CI(n22265), .I0(n2849[22]), .I1(GND_net), .CO(n22266));
    SB_LUT4 Mux_102_i1_3_lut (.I0(ootx_payloads_0_173), .I1(ootx_payloads_1_173), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[173]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_102_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1339_14_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n22541), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1741_2 (.CI(VCC_net), .I0(n2851[7]), .I1(n25187), 
            .CO(n22653));
    SB_LUT4 add_154_23_lut (.I0(GND_net), .I1(n2849[21]), .I2(GND_net), 
            .I3(n22264), .O(n2851[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_298 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n75), .O(n588));
    defparam i1_2_lut_3_lut_4_lut_adj_298.LUT_INIT = 16'h0100;
    SB_LUT4 i7132_3_lut_4_lut (.I0(n964), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_221), .O(n11242));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7132_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_736_8_lut (.I0(n1007), .I1(n1007), .I2(n1037), 
            .I3(n22418), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_14 (.CI(n22541), .I0(n1901), .I1(n1928), 
            .CO(n22542));
    SB_LUT4 mod_155_add_1674_25_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n22652), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_299 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n77), .O(n590));
    defparam i1_2_lut_3_lut_4_lut_adj_299.LUT_INIT = 16'h0100;
    SB_LUT4 Mux_103_i1_3_lut (.I0(ootx_payloads_0_172), .I1(ootx_payloads_1_172), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[172]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_103_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_104_i1_3_lut (.I0(ootx_payloads_0_171), .I1(ootx_payloads_1_171), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[171]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_104_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_105_i1_3_lut (.I0(ootx_payloads_0_170), .I1(ootx_payloads_1_170), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[170]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_105_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1339_13_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n22540), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_736_8 (.CI(n22418), .I0(n1007), .I1(n1037), .CO(n22419));
    SB_CARRY add_154_23 (.CI(n22264), .I0(n2849[21]), .I1(GND_net), .CO(n22265));
    SB_LUT4 Mux_106_i1_3_lut (.I0(ootx_payloads_0_169), .I1(ootx_payloads_1_169), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[169]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_106_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_107_i1_3_lut (.I0(ootx_payloads_0_168), .I1(ootx_payloads_1_168), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[168]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_107_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_736_7_lut (.I0(n1008_c), .I1(n1008_c), .I2(n1037), 
            .I3(n22417), .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_13 (.CI(n22540), .I0(n1902), .I1(n1928), 
            .CO(n22541));
    SB_LUT4 i1_2_lut_3_lut_adj_300 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n218), .I3(GND_net), .O(n602));
    defparam i1_2_lut_3_lut_adj_300.LUT_INIT = 16'h1010;
    SB_LUT4 EnabledDecoder_2_i58_2_lut_3_lut (.I0(n18_adj_1865), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n58_adj_2048));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i58_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_CARRY mod_155_add_1875_25 (.CI(n22724), .I0(n2690), .I1(n2720), 
            .CO(n22725));
    SB_CARRY mod_155_add_736_7 (.CI(n22417), .I0(n1008_c), .I1(n1037), 
            .CO(n22418));
    SB_LUT4 mod_155_add_1875_24_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n22723), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_108_i1_3_lut (.I0(ootx_payloads_0_167), .I1(ootx_payloads_1_167), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[167]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_108_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_301 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n220), .I3(GND_net), .O(n604));
    defparam i1_2_lut_3_lut_adj_301.LUT_INIT = 16'h1010;
    SB_LUT4 EnabledDecoder_2_i57_2_lut_3_lut (.I0(n18_adj_1865), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n57_adj_2045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i57_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mod_155_add_1674_24_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n22651), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_24 (.CI(n22651), .I0(n2391), .I1(n2423), 
            .CO(n22652));
    SB_LUT4 mod_155_add_1674_23_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n22650), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_adj_302 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n226), .I3(GND_net), .O(n610));
    defparam i1_2_lut_3_lut_adj_302.LUT_INIT = 16'h1010;
    SB_LUT4 Mux_109_i1_3_lut (.I0(ootx_payloads_0_166), .I1(ootx_payloads_1_166), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[166]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_109_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_110_i1_3_lut (.I0(ootx_payloads_0_165), .I1(ootx_payloads_1_165), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[165]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_110_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1339_12_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n22539), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_12 (.CI(n22539), .I0(n1903), .I1(n1928), 
            .CO(n22540));
    SB_LUT4 mod_155_add_736_6_lut (.I0(n1009), .I1(n1009), .I2(n25193), 
            .I3(n22416), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_736_6 (.CI(n22416), .I0(n1009), .I1(n25193), 
            .CO(n22417));
    SB_LUT4 i7723_3_lut_4_lut (.I0(n962), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1213), .O(n11833));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7723_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7131_3_lut_4_lut (.I0(n962), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_220), .O(n11241));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7131_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1339_11_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n22538), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_11 (.CI(n22538), .I0(n1904), .I1(n1928), 
            .CO(n22539));
    SB_LUT4 add_154_22_lut (.I0(GND_net), .I1(n2849[20]), .I2(GND_net), 
            .I3(n22263), .O(n2851[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 PrioSelect_33_i2_3_lut (.I0(data), .I1(n4485[3]), .I2(n34[0]), 
            .I3(GND_net), .O(n66_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_33_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_111_i1_3_lut (.I0(ootx_payloads_0_164), .I1(ootx_payloads_1_164), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[164]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_111_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_736_5_lut (.I0(n1010_c), .I1(n1010_c), .I2(n1037), 
            .I3(n22415), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_736_5 (.CI(n22415), .I0(n1010_c), .I1(n1037), 
            .CO(n22416));
    SB_CARRY add_66_23 (.CI(n22234), .I0(ootx_payloads_N_1699[21]), .I1(GND_net), 
            .CO(n22235));
    SB_LUT4 i1_2_lut_3_lut_adj_303 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n234), .I3(GND_net), .O(n618));
    defparam i1_2_lut_3_lut_adj_303.LUT_INIT = 16'h1010;
    SB_LUT4 i7118_3_lut_4_lut (.I0(n936), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_207), .O(n11228));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7118_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1674_23 (.CI(n22650), .I0(n2392), .I1(n2423), 
            .CO(n22651));
    SB_CARRY mod_155_add_2009_12 (.CI(n22764), .I0(n2903), .I1(n2918), 
            .CO(n22765));
    SB_LUT4 mod_155_add_1339_10_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n22537), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_112_i1_3_lut (.I0(ootx_payloads_0_163), .I1(ootx_payloads_1_163), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[163]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_112_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_113_i1_3_lut (.I0(ootx_payloads_0_162), .I1(ootx_payloads_1_162), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[162]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_113_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_736_4_lut (.I0(n1011), .I1(n1011), .I2(n1037), 
            .I3(n22414), .O(n1110)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_24 (.CI(n22723), .I0(n2691), .I1(n2720), 
            .CO(n22724));
    SB_LUT4 add_66_22_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[20]), 
            .I2(GND_net), .I3(n22233), .O(n337[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2009_11_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n22763), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7565_3_lut_4_lut (.I0(n646), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1371), .O(n11675));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1339_10 (.CI(n22537), .I0(n1905), .I1(n1928), 
            .CO(n22538));
    SB_LUT4 mod_155_add_1674_22_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n22649), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_154_22 (.CI(n22263), .I0(n2849[20]), .I1(GND_net), .CO(n22264));
    SB_LUT4 Mux_114_i1_3_lut (.I0(ootx_payloads_0_161), .I1(ootx_payloads_1_161), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[161]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_114_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_115_i1_3_lut (.I0(ootx_payloads_0_160), .I1(ootx_payloads_1_160), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[160]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_115_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_736_4 (.CI(n22414), .I0(n1011), .I1(n1037), .CO(n22415));
    SB_LUT4 mod_155_add_1339_9_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n22536), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_adj_304 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n250), .I3(GND_net), .O(n634));
    defparam i1_2_lut_3_lut_adj_304.LUT_INIT = 16'h1010;
    SB_CARRY mod_155_add_2143_24 (.CI(n22833), .I0(n3092), .I1(n3116), 
            .CO(n22834));
    SB_LUT4 mod_155_add_736_3_lut (.I0(n1012_c), .I1(n1012_c), .I2(n1037), 
            .I3(n22413), .O(n1111)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_3_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_66_22 (.CI(n22233), .I0(ootx_payloads_N_1699[20]), .I1(GND_net), 
            .CO(n22234));
    SB_LUT4 i1_2_lut_3_lut_adj_305 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n252), .I3(GND_net), .O(n636));
    defparam i1_2_lut_3_lut_adj_305.LUT_INIT = 16'h1010;
    SB_CARRY mod_155_add_2076_17 (.CI(n22797), .I0(n2998), .I1(n3017), 
            .CO(n22798));
    SB_CARRY mod_155_add_1339_9 (.CI(n22536), .I0(n1906), .I1(n1928), 
            .CO(n22537));
    SB_CARRY add_66_7 (.CI(n22218), .I0(\ootx_payloads_N_1699[5] ), .I1(GND_net), 
            .CO(n22219));
    SB_LUT4 i1_2_lut_3_lut_adj_306 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n256), .I3(GND_net), .O(n640));
    defparam i1_2_lut_3_lut_adj_306.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_307 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n79), .O(n720));
    defparam i1_2_lut_3_lut_4_lut_adj_307.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_116_i1_3_lut (.I0(ootx_payloads_0_159), .I1(ootx_payloads_1_159), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[159]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_116_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2009_11 (.CI(n22763), .I0(n2904), .I1(n2918), 
            .CO(n22764));
    SB_LUT4 i7030_3_lut_4_lut (.I0(n760), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_119), .O(n11140));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7030_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1875_23_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n22722), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_736_3 (.CI(n22413), .I0(n1012_c), .I1(n1037), 
            .CO(n22414));
    SB_LUT4 Mux_117_i1_3_lut (.I0(ootx_payloads_0_158), .I1(ootx_payloads_1_158), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[158]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_117_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7622_3_lut_4_lut (.I0(n760), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1314), .O(n11732));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7622_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1674_22 (.CI(n22649), .I0(n2393), .I1(n2423), 
            .CO(n22650));
    SB_LUT4 mod_155_add_1674_21_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n22648), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_2_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n337[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_308 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n258), .I3(GND_net), .O(n642));
    defparam i1_2_lut_3_lut_adj_308.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_309 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n260), .I3(GND_net), .O(n644));
    defparam i1_2_lut_3_lut_adj_309.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_310 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n262), .I3(GND_net), .O(n646));
    defparam i1_2_lut_3_lut_adj_310.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1339_8_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n22535), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_8 (.CI(n22535), .I0(n1907), .I1(n1928), 
            .CO(n22536));
    SB_LUT4 add_66_5_lut (.I0(GND_net), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(GND_net), .I3(n22216), .O(n337[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_736_2_lut (.I0(n2851[22]), .I1(n2851[22]), .I2(n25193), 
            .I3(VCC_net), .O(n1112)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_736_2 (.CI(VCC_net), .I0(n2851[22]), .I1(n25193), 
            .CO(n22413));
    SB_CARRY add_66_2 (.CI(VCC_net), .I0(ootx_payloads_N_1699[0]), .I1(GND_net), 
            .CO(n22214));
    SB_LUT4 Mux_118_i1_3_lut (.I0(ootx_payloads_0_157), .I1(ootx_payloads_1_157), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[157]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_118_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1339_7_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n22534), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1339_7 (.CI(n22534), .I0(n1908), .I1(n1928), 
            .CO(n22535));
    SB_CARRY add_66_6 (.CI(n22217), .I0(\ootx_payloads_N_1699[4] ), .I1(GND_net), 
            .CO(n22218));
    SB_LUT4 Mux_119_i1_3_lut (.I0(ootx_payloads_0_156), .I1(ootx_payloads_1_156), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[156]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_119_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_120_i1_3_lut (.I0(ootx_payloads_0_155), .I1(ootx_payloads_1_155), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[155]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_120_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_121_i1_3_lut (.I0(ootx_payloads_0_154), .I1(ootx_payloads_1_154), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[154]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_121_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_669_10_lut (.I0(n905), .I1(n905), .I2(n938_c), 
            .I3(n22412), .O(n1004_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_669_9_lut (.I0(n906_c), .I1(n906_c), .I2(n938_c), 
            .I3(n22411), .O(n1005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_122_i1_3_lut (.I0(ootx_payloads_0_153), .I1(ootx_payloads_1_153), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[153]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_122_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1674_21 (.CI(n22648), .I0(n2394), .I1(n2423), 
            .CO(n22649));
    SB_CARRY mod_155_add_1875_23 (.CI(n22722), .I0(n2692), .I1(n2720), 
            .CO(n22723));
    SB_LUT4 Mux_123_i1_3_lut (.I0(ootx_payloads_0_152), .I1(ootx_payloads_1_152), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[152]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_123_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1339_6_lut (.I0(n1909), .I1(n1909), .I2(n25191), 
            .I3(n22533), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1674_20_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n22647), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_66_4_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[2]), .I2(GND_net), 
            .I3(n22215), .O(n337[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20312_4_lut (.I0(counter_from_last_rise[1]), .I1(n291), .I2(counter_from_last_rise[3]), 
            .I3(counter_from_last_rise[2]), .O(n24676));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i20312_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 EnabledDecoder_2_i120_2_lut_3_lut (.I0(n40_adj_2049), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n120));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i120_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 Mux_124_i1_3_lut (.I0(ootx_payloads_0_151), .I1(ootx_payloads_1_151), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[151]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_124_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_669_9 (.CI(n22411), .I0(n906_c), .I1(n938_c), 
            .CO(n22412));
    SB_CARRY mod_155_add_1339_6 (.CI(n22533), .I0(n1909), .I1(n25191), 
            .CO(n22534));
    SB_LUT4 mod_155_add_1339_5_lut (.I0(n1910), .I1(n1910), .I2(n1928), 
            .I3(n22532), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_669_8_lut (.I0(n907), .I1(n907), .I2(n938_c), 
            .I3(n22410), .O(n1006_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_125_i1_3_lut (.I0(ootx_payloads_0_150), .I1(ootx_payloads_1_150), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[150]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_125_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i119_2_lut_3_lut (.I0(n40_adj_2049), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i119_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY mod_155_add_669_8 (.CI(n22410), .I0(n907), .I1(n938_c), .CO(n22411));
    SB_CARRY mod_155_add_1339_5 (.CI(n22532), .I0(n1910), .I1(n1928), 
            .CO(n22533));
    SB_LUT4 add_66_21_lut (.I0(GND_net), .I1(ootx_payloads_N_1699[19]), 
            .I2(GND_net), .I3(n22232), .O(n337[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_66_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1875_22_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n22721), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_669_7_lut (.I0(n908_c), .I1(n908_c), .I2(n938_c), 
            .I3(n22409), .O(n1007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_20 (.CI(n22647), .I0(n2395), .I1(n2423), 
            .CO(n22648));
    SB_LUT4 i1_2_lut_3_lut_adj_311 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n161), .I3(GND_net), .O(n674));
    defparam i1_2_lut_3_lut_adj_311.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_312 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n163), .I3(GND_net), .O(n676));
    defparam i1_2_lut_3_lut_adj_312.LUT_INIT = 16'h1010;
    SB_LUT4 Mux_126_i1_3_lut (.I0(ootx_payloads_0_149), .I1(ootx_payloads_1_149), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[149]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_126_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1674_19_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n22646), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_19 (.CI(n22646), .I0(n2396), .I1(n2423), 
            .CO(n22647));
    SB_LUT4 Mux_127_i1_3_lut (.I0(ootx_payloads_0_148), .I1(ootx_payloads_1_148), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[148]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_127_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1339_4_lut (.I0(n1911), .I1(n1911), .I2(n1928), 
            .I3(n22531), .O(n2010)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13599_4_lut (.I0(n24682), .I1(\counter_from_last_rise[8] ), 
            .I2(\counter_from_last_rise[6] ), .I3(counter_from_last_rise[4]), 
            .O(n119_adj_2050));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i13599_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 Mux_128_i1_3_lut (.I0(ootx_payloads_0_147), .I1(ootx_payloads_1_147), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[147]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_128_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7722_3_lut_4_lut (.I0(n960), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1214), .O(n11832));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7722_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_129_i1_3_lut (.I0(ootx_payloads_0_146), .I1(ootx_payloads_1_146), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[146]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_129_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_669_7 (.CI(n22409), .I0(n908_c), .I1(n938_c), 
            .CO(n22410));
    SB_CARRY mod_155_add_1339_4 (.CI(n22531), .I0(n1911), .I1(n1928), 
            .CO(n22532));
    SB_LUT4 add_154_21_lut (.I0(GND_net), .I1(n2849[19]), .I2(GND_net), 
            .I3(n22262), .O(n2851[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_154_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_313 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n165), .I3(GND_net), .O(n678));
    defparam i1_2_lut_3_lut_adj_313.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1339_3_lut (.I0(n1912), .I1(n1912), .I2(n1928), 
            .I3(n22530), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_669_6_lut (.I0(n909), .I1(n909), .I2(n25195), 
            .I3(n22408), .O(n1008_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_66_21 (.CI(n22232), .I0(ootx_payloads_N_1699[19]), .I1(GND_net), 
            .CO(n22233));
    SB_LUT4 i1_4_lut_adj_314 (.I0(n193_adj_2051), .I1(\counter_from_last_rise[11] ), 
            .I2(\counter_from_last_rise[8] ), .I3(\counter_from_last_rise[7] ), 
            .O(n4_adj_2052));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(251[8] 328[15])
    defparam i1_4_lut_adj_314.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_315 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n257), .I3(GND_net), .O(n770));
    defparam i1_2_lut_3_lut_adj_315.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_316 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n259), .I3(GND_net), .O(n772));
    defparam i1_2_lut_3_lut_adj_316.LUT_INIT = 16'h1010;
    SB_LUT4 i7130_3_lut_4_lut (.I0(n960), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_219), .O(n11240));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7130_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_130_i1_3_lut (.I0(ootx_payloads_0_145), .I1(ootx_payloads_1_145), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[145]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_130_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_317 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n261), .I3(GND_net), .O(n774));
    defparam i1_2_lut_3_lut_adj_317.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_318 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n77), .O(n718));
    defparam i1_2_lut_3_lut_4_lut_adj_318.LUT_INIT = 16'h1000;
    SB_CARRY mod_155_add_669_6 (.CI(n22408), .I0(n909), .I1(n25195), .CO(n22409));
    SB_CARRY mod_155_add_1339_3 (.CI(n22530), .I0(n1912), .I1(n1928), 
            .CO(n22531));
    SB_LUT4 i242_4_lut (.I0(\counter_from_last_rise[6] ), .I1(\counter_from_last_rise[7] ), 
            .I2(counter_from_last_rise[4]), .I3(counter_from_last_rise_c[5]), 
            .O(n283));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i242_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_319 (.I0(\counter_from_last_rise[9] ), .I1(\counter_from_last_rise[10] ), 
            .I2(n223), .I3(GND_net), .O(n256_adj_2053));
    defparam i1_3_lut_adj_319.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_320 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n167), .I3(GND_net), .O(n680));
    defparam i1_2_lut_3_lut_adj_320.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1674_18_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n22645), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_669_5_lut (.I0(n910_c), .I1(n910_c), .I2(n938_c), 
            .I3(n22407), .O(n1009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_131_i1_3_lut (.I0(ootx_payloads_0_144), .I1(ootx_payloads_1_144), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[144]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_131_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_132_i1_3_lut (.I0(ootx_payloads_0_143), .I1(ootx_payloads_1_143), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[143]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_132_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7575_3_lut_4_lut (.I0(n666), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1361), .O(n11685));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_321 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n169), .I3(GND_net), .O(n682));
    defparam i1_2_lut_3_lut_adj_321.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_322 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n171), .I3(GND_net), .O(n684));
    defparam i1_2_lut_3_lut_adj_322.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1339_2_lut (.I0(n2851[13]), .I1(n2851[13]), .I2(n25191), 
            .I3(VCC_net), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_2076_16_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n22796), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 PrioSelect_29_i2_3_lut (.I0(data), .I1(n4485[2]), .I2(n34[0]), 
            .I3(GND_net), .O(n62_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_323 (.I0(\counter_from_last_rise[10] ), .I1(n283), 
            .I2(\counter_from_last_rise[9] ), .I3(\counter_from_last_rise[8] ), 
            .O(n24004));
    defparam i2_4_lut_adj_323.LUT_INIT = 16'h8000;
    SB_LUT4 Mux_133_i1_3_lut (.I0(ootx_payloads_0_142), .I1(ootx_payloads_1_142), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[142]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_133_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_324 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n112_adj_2043), .O(n688));
    defparam i1_2_lut_3_lut_4_lut_adj_324.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_325 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n116), .O(n564));
    defparam i1_2_lut_3_lut_4_lut_adj_325.LUT_INIT = 16'h0100;
    SB_LUT4 Mux_134_i1_3_lut (.I0(ootx_payloads_0_141), .I1(ootx_payloads_1_141), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[141]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_134_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_669_5 (.CI(n22407), .I0(n910_c), .I1(n938_c), 
            .CO(n22408));
    SB_LUT4 Mux_135_i1_3_lut (.I0(ootx_payloads_0_140), .I1(ootx_payloads_1_140), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[140]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_135_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_326 (.I0(ootx_payloads_N_1699[0]), .I1(n8941), 
            .I2(n88), .I3(GND_net), .O(n6_adj_2054));
    defparam i1_3_lut_adj_326.LUT_INIT = 16'h0202;
    SB_CARRY mod_155_add_1339_2 (.CI(VCC_net), .I0(n2851[13]), .I1(n25191), 
            .CO(n22530));
    SB_LUT4 mod_155_add_2009_10_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n22762), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut_adj_327 (.I0(\counter_from_last_rise[10] ), .I1(\counter_from_last_rise[12] ), 
            .I2(n4_adj_2052), .I3(\counter_from_last_rise[9] ), .O(n7));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(251[8] 328[15])
    defparam i1_4_lut_adj_327.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_328 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n118_adj_2055), .O(n566));
    defparam i1_2_lut_3_lut_4_lut_adj_328.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_329 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n118_adj_2055), .O(n694));
    defparam i1_2_lut_3_lut_4_lut_adj_329.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_330 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n120), .O(n568));
    defparam i1_2_lut_3_lut_4_lut_adj_330.LUT_INIT = 16'h0100;
    SB_LUT4 mod_155_add_669_4_lut (.I0(n911), .I1(n911), .I2(n938_c), 
            .I3(n22406), .O(n1010_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_22 (.CI(n22721), .I0(n2693), .I1(n2720), 
            .CO(n22722));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_331 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n122_adj_2046), .O(n570));
    defparam i1_2_lut_3_lut_4_lut_adj_331.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_332 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n124), .O(n572));
    defparam i1_2_lut_3_lut_4_lut_adj_332.LUT_INIT = 16'h0100;
    SB_CARRY mod_155_add_2009_10 (.CI(n22762), .I0(n2905), .I1(n2918), 
            .CO(n22763));
    SB_CARRY mod_155_add_1674_18 (.CI(n22645), .I0(n2397), .I1(n2423), 
            .CO(n22646));
    SB_LUT4 i1_4_lut_adj_333 (.I0(\counter_from_last_rise[12] ), .I1(\counter_from_last_rise[11] ), 
            .I2(n24004), .I3(n256_adj_2053), .O(n5));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(251[8] 328[15])
    defparam i1_4_lut_adj_333.LUT_INIT = 16'ha888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_334 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n126_adj_1853), .O(n574));
    defparam i1_2_lut_3_lut_4_lut_adj_334.LUT_INIT = 16'h0100;
    SB_LUT4 i6983_3_lut_4_lut (.I0(n666), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_72), .O(n11093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1875_21_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n22720), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1272_19_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n22529), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_i405_3_lut_4_lut (.I0(n19313), .I1(n83), .I2(n58_adj_1820), 
            .I3(n2851[29]), .O(n610_c));
    defparam mod_155_i405_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 i1_4_lut_adj_335 (.I0(n9029), .I1(n5), .I2(n19257), .I3(n7), 
            .O(data_N_1765));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(251[8] 328[15])
    defparam i1_4_lut_adj_335.LUT_INIT = 16'hefee;
    SB_LUT4 Mux_136_i1_3_lut (.I0(ootx_payloads_0_139), .I1(ootx_payloads_1_139), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[139]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_136_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_i406_3_lut_4_lut (.I0(n19313), .I1(n83), .I2(n2851[27]), 
            .I3(n2851[28]), .O(n611));
    defparam mod_155_i406_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 mod_155_add_1674_17_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n22644), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_669_4 (.CI(n22406), .I0(n911), .I1(n938_c), .CO(n22407));
    SB_LUT4 Mux_137_i1_3_lut (.I0(ootx_payloads_0_138), .I1(ootx_payloads_1_138), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[138]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_137_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_336 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n132), .O(n580));
    defparam i1_2_lut_3_lut_4_lut_adj_336.LUT_INIT = 16'h0100;
    SB_LUT4 mod_155_i404_3_lut_4_lut (.I0(n19313), .I1(n83), .I2(n60_c), 
            .I3(n2851[30]), .O(n609));
    defparam mod_155_i404_3_lut_4_lut.LUT_INIT = 16'hf708;
    SB_LUT4 Mux_138_i1_3_lut (.I0(ootx_payloads_0_137), .I1(ootx_payloads_1_137), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[137]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_138_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_337 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n134_adj_1948), .O(n582));
    defparam i1_2_lut_3_lut_4_lut_adj_337.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_338 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n73), .O(n586));
    defparam i1_2_lut_3_lut_4_lut_adj_338.LUT_INIT = 16'h0100;
    SB_LUT4 Mux_139_i1_3_lut (.I0(ootx_payloads_0_136), .I1(ootx_payloads_1_136), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[136]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_139_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 PrioSelect_25_i2_3_lut (.I0(data), .I1(n4485[1]), .I2(n34[0]), 
            .I3(GND_net), .O(n58_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_25_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_339 (.I0(n19313), .I1(n83), .I2(n2851[27]), 
            .I3(GND_net), .O(n612_c));
    defparam i1_2_lut_3_lut_adj_339.LUT_INIT = 16'h7878;
    SB_LUT4 Mux_140_i1_3_lut (.I0(ootx_payloads_0_135), .I1(ootx_payloads_1_135), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[135]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_140_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1272_18_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n22528), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1272_18 (.CI(n22528), .I0(n1797), .I1(n1829), 
            .CO(n22529));
    SB_LUT4 mod_155_add_669_3_lut (.I0(n912_c), .I1(n912_c), .I2(n938_c), 
            .I3(n22405), .O(n1011)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_3_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_669_3 (.CI(n22405), .I0(n912_c), .I1(n938_c), 
            .CO(n22406));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_340 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n125), .O(n766));
    defparam i1_2_lut_3_lut_4_lut_adj_340.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_1272_17_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n22527), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_17 (.CI(n22644), .I0(n2398), .I1(n2423), 
            .CO(n22645));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_341 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n93_adj_2014), .O(n734));
    defparam i1_2_lut_3_lut_4_lut_adj_341.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_342 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n135), .O(n776));
    defparam i1_2_lut_3_lut_4_lut_adj_342.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_141_i1_3_lut (.I0(ootx_payloads_0_134), .I1(ootx_payloads_1_134), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[134]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_141_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_142_i1_3_lut (.I0(ootx_payloads_0_133), .I1(ootx_payloads_1_133), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[133]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_142_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_143_i1_3_lut (.I0(ootx_payloads_0_132), .I1(ootx_payloads_1_132), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[132]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_143_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_144_i1_3_lut (.I0(ootx_payloads_0_131), .I1(ootx_payloads_1_131), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[131]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_144_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_669_2_lut (.I0(n2851[23]), .I1(n2851[23]), .I2(n25195), 
            .I3(VCC_net), .O(n1012_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_669_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1272_17 (.CI(n22527), .I0(n1798), .I1(n1829), 
            .CO(n22528));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_343 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n90_adj_1876), .O(n538));
    defparam i1_2_lut_3_lut_4_lut_adj_343.LUT_INIT = 16'h0100;
    SB_LUT4 mod_155_add_1674_16_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n22643), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_669_2 (.CI(VCC_net), .I0(n2851[23]), .I1(n25195), 
            .CO(n22405));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_344 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n115), .O(n756));
    defparam i1_2_lut_3_lut_4_lut_adj_344.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_345 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n117), .O(n758));
    defparam i1_2_lut_3_lut_4_lut_adj_345.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_145_i1_3_lut (.I0(ootx_payloads_0_130), .I1(ootx_payloads_1_130), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[130]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_145_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1272_16_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n22526), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1272_16 (.CI(n22526), .I0(n1799), .I1(n1829), 
            .CO(n22527));
    SB_LUT4 Mux_146_i1_3_lut (.I0(ootx_payloads_0_129), .I1(ootx_payloads_1_129), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[129]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_146_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_346 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n136), .O(n712));
    defparam i1_2_lut_3_lut_4_lut_adj_346.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_602_9_lut (.I0(GND_net), .I1(n806_c), .I2(VCC_net), 
            .I3(n22404), .O(n71[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_602_8_lut (.I0(GND_net), .I1(n807), .I2(VCC_net), 
            .I3(n22403), .O(n71[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut (.I0(n36_adj_2041), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n84));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i84_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_347 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n87), .O(n728));
    defparam i1_2_lut_3_lut_4_lut_adj_347.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_147_i1_3_lut (.I0(ootx_payloads_0_128), .I1(ootx_payloads_1_128), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[128]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_147_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1272_15_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n22525), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_21 (.CI(n22720), .I0(n2694), .I1(n2720), 
            .CO(n22721));
    SB_LUT4 Mux_148_i1_3_lut (.I0(ootx_payloads_0_127), .I1(ootx_payloads_1_127), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[127]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_148_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_348 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n73), .O(n714));
    defparam i1_2_lut_3_lut_4_lut_adj_348.LUT_INIT = 16'h1000;
    SB_CARRY mod_155_add_602_8 (.CI(n22403), .I0(n807), .I1(VCC_net), 
            .CO(n22404));
    SB_LUT4 i1_2_lut_3_lut_adj_349 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n217), .I3(GND_net), .O(n730));
    defparam i1_2_lut_3_lut_adj_349.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1875_20_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n22719), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_16 (.CI(n22643), .I0(n2399), .I1(n2423), 
            .CO(n22644));
    SB_LUT4 EnabledDecoder_3_i2_2_lut (.I0(n432), .I1(\lighthouse[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n34[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(126[25:35])
    defparam EnabledDecoder_3_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_350 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n219), .I3(GND_net), .O(n732));
    defparam i1_2_lut_3_lut_adj_350.LUT_INIT = 16'h1010;
    SB_LUT4 Mux_149_i1_3_lut (.I0(ootx_payloads_0_126), .I1(ootx_payloads_1_126), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[126]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_149_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1674_15_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n22642), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1272_15 (.CI(n22525), .I0(n1800), .I1(n1829), 
            .CO(n22526));
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut (.I0(n36_adj_2041), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n83_adj_2035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i83_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 Mux_150_i1_3_lut (.I0(ootx_payloads_0_125), .I1(ootx_payloads_1_125), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[125]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_150_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1272_14_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n22524), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_602_7_lut (.I0(GND_net), .I1(n808_c), .I2(VCC_net), 
            .I3(n22402), .O(n71[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Mux_151_i1_3_lut (.I0(ootx_payloads_0_124), .I1(ootx_payloads_1_124), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[124]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_151_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_152_i1_3_lut (.I0(ootx_payloads_0_123), .I1(ootx_payloads_1_123), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[123]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_152_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_153_i1_3_lut (.I0(ootx_payloads_0_122), .I1(ootx_payloads_1_122), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[122]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_153_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_602_7 (.CI(n22402), .I0(n808_c), .I1(VCC_net), 
            .CO(n22403));
    SB_CARRY mod_155_add_1272_14 (.CI(n22524), .I0(n1801), .I1(n1829), 
            .CO(n22525));
    SB_LUT4 EnabledDecoder_3_i3_2_lut (.I0(n432), .I1(\lighthouse[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n34[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(126[25:35])
    defparam EnabledDecoder_3_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_351 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n75), .O(n716));
    defparam i1_2_lut_3_lut_4_lut_adj_351.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_1272_13_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n22523), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_602_6_lut (.I0(GND_net), .I1(n809), .I2(GND_net), 
            .I3(n22401), .O(n71[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_352 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n114_adj_2044), .O(n562));
    defparam i1_2_lut_3_lut_4_lut_adj_352.LUT_INIT = 16'h0100;
    SB_CARRY mod_155_add_602_6 (.CI(n22401), .I0(n809), .I1(GND_net), 
            .CO(n22402));
    SB_LUT4 i1_2_lut_3_lut_adj_353 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n225), .I3(GND_net), .O(n738));
    defparam i1_2_lut_3_lut_adj_353.LUT_INIT = 16'h1010;
    SB_CARRY mod_155_add_1674_15 (.CI(n22642), .I0(n2400), .I1(n2423), 
            .CO(n22643));
    SB_LUT4 mod_155_add_1674_14_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n22641), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_154_i1_3_lut (.I0(ootx_payloads_0_121), .I1(ootx_payloads_1_121), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[121]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_154_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1272_13 (.CI(n22523), .I0(n1802), .I1(n1829), 
            .CO(n22524));
    SB_LUT4 mod_155_add_1272_12_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n22522), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7029_3_lut_4_lut (.I0(n758), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_118), .O(n11139));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7029_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_155_i1_3_lut (.I0(ootx_payloads_0_120), .I1(ootx_payloads_1_120), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[120]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_155_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_602_5_lut (.I0(GND_net), .I1(n810_c), .I2(VCC_net), 
            .I3(n22400), .O(n71[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_602_5 (.CI(n22400), .I0(n810_c), .I1(VCC_net), 
            .CO(n22401));
    SB_LUT4 Mux_156_i1_3_lut (.I0(ootx_payloads_0_119), .I1(ootx_payloads_1_119), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[119]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_156_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1272_12 (.CI(n22522), .I0(n1803), .I1(n1829), 
            .CO(n22523));
    SB_LUT4 mod_155_add_1272_11_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n22521), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_157_i1_3_lut (.I0(ootx_payloads_0_118), .I1(ootx_payloads_1_118), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[118]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_157_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_602_4_lut (.I0(GND_net), .I1(n811), .I2(VCC_net), 
            .I3(n22399), .O(n71[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_602_4 (.CI(n22399), .I0(n811), .I1(VCC_net), 
            .CO(n22400));
    SB_LUT4 Mux_158_i1_3_lut (.I0(ootx_payloads_0_117), .I1(ootx_payloads_1_117), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[117]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_158_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_354 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n233), .I3(GND_net), .O(n746));
    defparam i1_2_lut_3_lut_adj_354.LUT_INIT = 16'h1010;
    SB_LUT4 Mux_159_i1_3_lut (.I0(ootx_payloads_0_116), .I1(ootx_payloads_1_116), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[116]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_159_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20469_2_lut (.I0(reset_c), .I1(new_data), .I2(GND_net), .I3(GND_net), 
            .O(n18844));
    defparam i20469_2_lut.LUT_INIT = 16'h1111;
    SB_CARRY mod_155_add_2076_16 (.CI(n22796), .I0(n2999), .I1(n3017), 
            .CO(n22797));
    SB_LUT4 mod_155_add_2009_9_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n22761), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_160_i1_3_lut (.I0(ootx_payloads_0_115), .I1(ootx_payloads_1_115), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[115]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_160_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7621_3_lut_4_lut (.I0(n758), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1315), .O(n11731));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7621_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2009_9 (.CI(n22761), .I0(n2906), .I1(n2918), 
            .CO(n22762));
    SB_CARRY mod_155_add_1875_20 (.CI(n22719), .I0(n2695), .I1(n2720), 
            .CO(n22720));
    SB_LUT4 Mux_161_i1_3_lut (.I0(ootx_payloads_0_114), .I1(ootx_payloads_1_114), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[114]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_161_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1875_19_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n22718), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_14 (.CI(n22641), .I0(n2401), .I1(n2423), 
            .CO(n22642));
    SB_LUT4 mod_155_add_2009_8_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n22760), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_355 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n81), .O(n722));
    defparam i1_2_lut_3_lut_4_lut_adj_355.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_162_i1_3_lut (.I0(ootx_payloads_0_113), .I1(ootx_payloads_1_113), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[113]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_162_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1674_13_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n22640), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1272_11 (.CI(n22521), .I0(n1804), .I1(n1829), 
            .CO(n22522));
    SB_LUT4 mod_155_add_1272_10_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n22520), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_602_3_lut (.I0(GND_net), .I1(n812_c), .I2(VCC_net), 
            .I3(n22398), .O(n71[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_356 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n119), .O(n760));
    defparam i1_2_lut_3_lut_4_lut_adj_356.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_163_i1_3_lut (.I0(ootx_payloads_0_112), .I1(ootx_payloads_1_112), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[112]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_163_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_602_3 (.CI(n22398), .I0(n812_c), .I1(VCC_net), 
            .CO(n22399));
    SB_CARRY mod_155_add_1272_10 (.CI(n22520), .I0(n1805), .I1(n1829), 
            .CO(n22521));
    SB_CARRY mod_155_add_2009_8 (.CI(n22760), .I0(n2907), .I1(n2918), 
            .CO(n22761));
    SB_LUT4 i7011_3_lut_4_lut (.I0(n722), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_100), .O(n11121));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7011_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_357 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n83_adj_2035), .O(n724));
    defparam i1_2_lut_3_lut_4_lut_adj_357.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_1272_9_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n22519), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_602_2_lut (.I0(GND_net), .I1(n2851[24]), .I2(GND_net), 
            .I3(VCC_net), .O(n71[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_602_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Mux_22_i1_3_lut_adj_358 (.I0(bit_counters_0_14), .I1(bit_counters_1_14), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[14]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_22_i1_3_lut_adj_358.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_359 (.I0(sensor_state_switch_counter[5]), .I1(n2276), 
            .I2(n37_adj_1914), .I3(sensor_state_switch_counter[3]), .O(n10_adj_2057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(199[5] 341[12])
    defparam i4_4_lut_adj_359.LUT_INIT = 16'hfffb;
    SB_LUT4 Mux_164_i1_3_lut (.I0(ootx_payloads_0_111), .I1(ootx_payloads_1_111), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[111]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_164_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7603_3_lut_4_lut (.I0(n722), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1333), .O(n11713));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7603_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_602_2 (.CI(VCC_net), .I0(n2851[24]), .I1(GND_net), 
            .CO(n22398));
    SB_CARRY mod_155_add_1674_13 (.CI(n22640), .I0(n2402), .I1(n2423), 
            .CO(n22641));
    SB_LUT4 i1_2_lut_3_lut_adj_360 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n249), .I3(GND_net), .O(n762));
    defparam i1_2_lut_3_lut_adj_360.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_361 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n251), .I3(GND_net), .O(n764));
    defparam i1_2_lut_3_lut_adj_361.LUT_INIT = 16'h1010;
    SB_LUT4 mod_155_add_1674_12_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n22639), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_165_i1_3_lut (.I0(ootx_payloads_0_110), .I1(ootx_payloads_1_110), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[110]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_165_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1272_9 (.CI(n22519), .I0(n1806), .I1(n1829), 
            .CO(n22520));
    SB_LUT4 mod_155_add_1272_8_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n22518), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2076_15_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n22795), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_362 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n85), .O(n726));
    defparam i1_2_lut_3_lut_4_lut_adj_362.LUT_INIT = 16'h1000;
    SB_LUT4 mod_155_add_535_8_lut (.I0(n740_c), .I1(n707), .I2(VCC_net), 
            .I3(n22397), .O(n806_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_155_add_535_7_lut (.I0(GND_net), .I1(n708_c), .I2(VCC_net), 
            .I3(n22396), .O(n773[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_2076_15 (.CI(n22795), .I0(n3000), .I1(n3017), 
            .CO(n22796));
    SB_LUT4 Mux_166_i1_3_lut (.I0(ootx_payloads_0_109), .I1(ootx_payloads_1_109), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[109]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_166_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_167_i1_3_lut (.I0(ootx_payloads_0_108), .I1(ootx_payloads_1_108), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[108]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_167_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_363 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n255), .I3(GND_net), .O(n768));
    defparam i1_2_lut_3_lut_adj_363.LUT_INIT = 16'h1010;
    SB_LUT4 Mux_168_i1_3_lut (.I0(ootx_payloads_0_107), .I1(ootx_payloads_1_107), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[107]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_168_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1272_8 (.CI(n22518), .I0(n1807), .I1(n1829), 
            .CO(n22519));
    SB_LUT4 mod_155_add_1272_7_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n22517), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20531_1_lut (.I0(n1631_adj_2058), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25199));
    defparam i20531_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i256_2_lut_3_lut (.I0(n63_adj_2059), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n256));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i256_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_CARRY mod_155_add_535_7 (.CI(n22396), .I0(n708_c), .I1(VCC_net), 
            .CO(n22397));
    SB_LUT4 mod_155_add_535_6_lut (.I0(GND_net), .I1(n709), .I2(GND_net), 
            .I3(n22395), .O(n773[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2143_23_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n22832), .O(n43_adj_1961)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i255_2_lut_3_lut (.I0(n63_adj_2059), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n255));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i255_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7518_3_lut_4_lut (.I0(n552), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1418), .O(n11628));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7518_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_169_i1_3_lut (.I0(ootx_payloads_0_106), .I1(ootx_payloads_1_106), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[106]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_169_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_170_i1_3_lut (.I0(ootx_payloads_0_105), .I1(ootx_payloads_1_105), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[105]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_170_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1875_19 (.CI(n22718), .I0(n2696), .I1(n2720), 
            .CO(n22719));
    SB_LUT4 mod_155_add_1875_18_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n22717), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_171_i1_3_lut (.I0(ootx_payloads_0_104), .I1(ootx_payloads_1_104), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[104]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_171_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1674_12 (.CI(n22639), .I0(n2403), .I1(n2423), 
            .CO(n22640));
    SB_CARRY mod_155_add_1272_7 (.CI(n22517), .I0(n1808), .I1(n1829), 
            .CO(n22518));
    SB_LUT4 mod_155_add_1674_11_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n22638), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6888_3_lut_4_lut (.I0(n552), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_15), .O(n10998));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i118_2_lut_3_lut (.I0(n38_c), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n118_adj_2055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i118_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 Mux_172_i1_3_lut (.I0(ootx_payloads_0_103), .I1(ootx_payloads_1_103), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[103]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_172_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_173_i1_3_lut (.I0(ootx_payloads_0_102), .I1(ootx_payloads_1_102), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[102]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_173_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_174_i1_3_lut (.I0(ootx_payloads_0_101), .I1(ootx_payloads_1_101), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[101]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_174_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_364 (.I0(n77), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n846));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_364.LUT_INIT = 16'h0020;
    SB_CARRY mod_155_add_535_6 (.CI(n22395), .I0(n709), .I1(GND_net), 
            .CO(n22396));
    SB_LUT4 mod_155_add_1272_6_lut (.I0(n1809), .I1(n1809), .I2(n25196), 
            .I3(n22516), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_155_add_1272_6 (.CI(n22516), .I0(n1809), .I1(n25196), 
            .CO(n22517));
    SB_LUT4 mod_155_add_535_5_lut (.I0(GND_net), .I1(n710_c), .I2(VCC_net), 
            .I3(n22394), .O(n773[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF i929_930 (.Q(n1216), .C(clock_c), .D(n11830));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_535_5 (.CI(n22394), .I0(n710_c), .I1(VCC_net), 
            .CO(n22395));
    SB_LUT4 mod_155_add_1272_5_lut (.I0(n1810), .I1(n1810), .I2(n1829), 
            .I3(n22515), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i117_2_lut_3_lut (.I0(n38_c), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i117_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY mod_155_add_1674_11 (.CI(n22638), .I0(n2404), .I1(n2423), 
            .CO(n22639));
    SB_LUT4 mod_155_add_535_4_lut (.I0(GND_net), .I1(n711), .I2(VCC_net), 
            .I3(n22393), .O(n773[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_2143_23 (.CI(n22832), .I0(n3093), .I1(n3116), 
            .CO(n22833));
    SB_LUT4 i7664_3_lut_4_lut (.I0(n844), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1272), .O(n11774));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7664_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i926_927 (.Q(n1217), .C(clock_c), .D(n11829));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_175_i1_3_lut (.I0(ootx_payloads_0_100), .I1(ootx_payloads_1_100), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[100]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_175_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1272_5 (.CI(n22515), .I0(n1810), .I1(n1829), 
            .CO(n22516));
    SB_LUT4 mod_155_add_1674_10_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n22637), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7072_3_lut_4_lut (.I0(n844), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_161), .O(n11182));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7072_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6973_3_lut_4_lut (.I0(n646), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_62), .O(n11083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i923_924 (.Q(n1218), .C(clock_c), .D(n11828));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_535_4 (.CI(n22393), .I0(n711), .I1(VCC_net), 
            .CO(n22394));
    SB_LUT4 mod_155_add_1272_4_lut (.I0(n1811), .I1(n1811), .I2(n1829), 
            .I3(n22514), .O(n1910)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2076_14_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n22794), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_176_i1_3_lut (.I0(ootx_payloads_0_99), .I1(ootx_payloads_1_99), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[99]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_176_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_365 (.I0(n75), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n844));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_365.LUT_INIT = 16'h0020;
    SB_CARRY mod_155_add_1272_4 (.CI(n22514), .I0(n1811), .I1(n1829), 
            .CO(n22515));
    SB_LUT4 mod_155_add_535_3_lut (.I0(GND_net), .I1(n712_c), .I2(VCC_net), 
            .I3(n22392), .O(n773[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2009_7_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n22759), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i920_921 (.Q(n1219), .C(clock_c), .D(n11827));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7663_3_lut_4_lut (.I0(n842), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1273), .O(n11773));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7663_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7071_3_lut_4_lut (.I0(n842), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_160), .O(n11181));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7071_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_535_3 (.CI(n22392), .I0(n712_c), .I1(VCC_net), 
            .CO(n22393));
    SB_LUT4 mod_155_add_1272_3_lut (.I0(n1812), .I1(n1812), .I2(n1829), 
            .I3(n22513), .O(n1911)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7517_3_lut_4_lut (.I0(n550), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1419), .O(n11627));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2009_7 (.CI(n22759), .I0(n2908), .I1(n2918), 
            .CO(n22760));
    SB_LUT4 mod_155_add_535_2_lut (.I0(GND_net), .I1(n2851[25]), .I2(GND_net), 
            .I3(VCC_net), .O(n773[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_535_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6889_3_lut_4_lut (.I0(n550), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_14), .O(n10999));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i917_918 (.Q(n1220), .C(clock_c), .D(n11826));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_177_i1_3_lut (.I0(ootx_payloads_0_98), .I1(ootx_payloads_1_98), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[98]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_177_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1875_18 (.CI(n22717), .I0(n2697), .I1(n2720), 
            .CO(n22718));
    SB_CARRY mod_155_add_2076_14 (.CI(n22794), .I0(n3001), .I1(n3017), 
            .CO(n22795));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_366 (.I0(n73), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n842));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_366.LUT_INIT = 16'h0020;
    SB_CARRY mod_155_add_1674_10 (.CI(n22637), .I0(n2405), .I1(n2423), 
            .CO(n22638));
    SB_LUT4 mod_155_add_2076_13_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n22793), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_178_i1_3_lut (.I0(ootx_payloads_0_97), .I1(ootx_payloads_1_97), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[97]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_178_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_179_i1_3_lut (.I0(ootx_payloads_0_96), .I1(ootx_payloads_1_96), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[96]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_179_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i914_915 (.Q(n1221), .C(clock_c), .D(n11825));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7003_3_lut_4_lut (.I0(n706), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_92), .O(n11113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7003_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1272_3 (.CI(n22513), .I0(n1812), .I1(n1829), 
            .CO(n22514));
    SB_LUT4 mod_155_add_2143_22_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n22831), .O(n41_adj_1959)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_180_i1_3_lut (.I0(ootx_payloads_0_95), .I1(ootx_payloads_1_95), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[95]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_180_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_535_2 (.CI(VCC_net), .I0(n2851[25]), .I1(GND_net), 
            .CO(n22392));
    SB_LUT4 Mux_181_i1_3_lut (.I0(ootx_payloads_0_94), .I1(ootx_payloads_1_94), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[94]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_181_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_182_i1_3_lut (.I0(ootx_payloads_0_93), .I1(ootx_payloads_1_93), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[93]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_182_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1272_2_lut (.I0(n2851[14]), .I1(n2851[14]), .I2(n25196), 
            .I3(VCC_net), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFF i911_912 (.Q(n1222), .C(clock_c), .D(n11824));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2076_13 (.CI(n22793), .I0(n3002), .I1(n3017), 
            .CO(n22794));
    SB_CARRY mod_155_add_2143_22 (.CI(n22831), .I0(n3094), .I1(n3116), 
            .CO(n22832));
    SB_LUT4 Mux_183_i1_3_lut (.I0(ootx_payloads_0_92), .I1(ootx_payloads_1_92), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[92]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_183_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_468_7_lut (.I0(n641), .I1(n608_c), .I2(VCC_net), 
            .I3(n22391), .O(n707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_468_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_155_add_2009_6_lut (.I0(n2909), .I1(n2909), .I2(n25182), 
            .I3(n22758), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i7595_3_lut_4_lut (.I0(n706), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1341), .O(n11705));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7595_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_184_i1_3_lut (.I0(ootx_payloads_0_91), .I1(ootx_payloads_1_91), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[91]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_184_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i908_909 (.Q(n1223), .C(clock_c), .D(n11823));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_185_i1_3_lut (.I0(ootx_payloads_0_90), .I1(ootx_payloads_1_90), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[90]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_185_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_367 (.I0(n130_adj_2047), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n962));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_367.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_1674_9_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n22636), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1875_17_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n22716), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1272_2 (.CI(VCC_net), .I0(n2851[14]), .I1(n25196), 
            .CO(n22513));
    SB_CARRY mod_155_add_1674_9 (.CI(n22636), .I0(n2406), .I1(n2423), 
            .CO(n22637));
    SB_DFF i905_906 (.Q(n1224), .C(clock_c), .D(n11822));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_468_6_lut (.I0(GND_net), .I1(n609), .I2(GND_net), 
            .I3(n22390), .O(n89[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_468_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_from_nskip_rise_640_add_4_7_lut (.I0(n6333_c[5]), .I1(n2280), 
            .I2(counter_from_nskip_rise[5]), .I3(n22355), .O(n91[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mod_155_add_2076_12_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n22792), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_186_i1_3_lut (.I0(ootx_payloads_0_89), .I1(ootx_payloads_1_89), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[89]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_186_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_187_i1_3_lut (.I0(ootx_payloads_0_88), .I1(ootx_payloads_1_88), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[88]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_187_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i37_2_lut_3_lut (.I0(n13_adj_1854), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(GND_net), .O(n37_adj_1949));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i37_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i902_903 (.Q(n1225), .C(clock_c), .D(n11821));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1205_18_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n22512), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_188_i1_3_lut (.I0(ootx_payloads_0_87), .I1(ootx_payloads_1_87), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[87]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_188_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_468_6 (.CI(n22390), .I0(n609), .I1(GND_net), 
            .CO(n22391));
    SB_CARRY counter_from_nskip_rise_640_add_4_7 (.CI(n22355), .I0(n2280), 
            .I1(counter_from_nskip_rise[5]), .CO(n22356));
    SB_LUT4 Mux_189_i1_3_lut (.I0(ootx_payloads_0_86), .I1(ootx_payloads_1_86), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[86]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_189_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7662_3_lut_4_lut (.I0(n840), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1274), .O(n11772));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7662_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_190_i1_3_lut (.I0(ootx_payloads_0_85), .I1(ootx_payloads_1_85), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[85]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_190_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1875_17 (.CI(n22716), .I0(n2698), .I1(n2720), 
            .CO(n22717));
    SB_LUT4 Mux_191_i1_3_lut (.I0(ootx_payloads_0_84), .I1(ootx_payloads_1_84), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[84]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_191_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i899_900 (.Q(n1226), .C(clock_c), .D(n11820));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_2143_21_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n22830), .O(n39_adj_1973)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7070_3_lut_4_lut (.I0(n840), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_159), .O(n11180));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7070_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_368 (.I0(n136), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n840));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_368.LUT_INIT = 16'h0020;
    SB_LUT4 mod_155_add_1674_8_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n22635), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_8 (.CI(n22635), .I0(n2407), .I1(n2423), 
            .CO(n22636));
    SB_LUT4 Mux_192_i1_3_lut (.I0(ootx_payloads_0_83), .I1(ootx_payloads_1_83), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[83]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_192_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7516_3_lut_4_lut (.I0(n548), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1420), .O(n11626));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7516_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_17_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n22511), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 counter_from_nskip_rise_640_add_4_6_lut (.I0(n6361), .I1(n2280), 
            .I2(counter_from_nskip_rise[4]), .I3(n22354), .O(n91[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_6_lut.LUT_INIT = 16'h8BB8;
    SB_DFF i896_897 (.Q(n1227), .C(clock_c), .D(n11819));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_468_5_lut (.I0(GND_net), .I1(n610_c), .I2(VCC_net), 
            .I3(n22389), .O(n89[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_468_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut (.I0(n13_adj_1854), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(GND_net), .O(n38_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i38_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i6891_3_lut_4_lut (.I0(n548), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_13), .O(n11001));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1875_16_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n22715), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_193_i1_3_lut (.I0(ootx_payloads_0_82), .I1(ootx_payloads_1_82), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[82]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_193_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i893_894 (.Q(n1228), .C(clock_c), .D(n11818));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7661_3_lut_4_lut (.I0(n838), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1275), .O(n11771));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7661_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_369 (.I0(ootx_payloads_N_1744[0]), .I1(n20105), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n72[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(188[20:30])
    defparam i2_3_lut_adj_369.LUT_INIT = 16'h8080;
    SB_LUT4 Mux_194_i1_3_lut (.I0(ootx_payloads_0_81), .I1(ootx_payloads_1_81), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[81]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_194_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1205_17 (.CI(n22511), .I0(n1698), .I1(n1730), 
            .CO(n22512));
    SB_CARRY counter_from_nskip_rise_640_add_4_6 (.CI(n22354), .I0(n2280), 
            .I1(counter_from_nskip_rise[4]), .CO(n22355));
    SB_LUT4 i7709_3_lut_4_lut (.I0(n934), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1227), .O(n11819));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7709_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7069_3_lut_4_lut (.I0(n838), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_158), .O(n11179));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7069_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_468_5 (.CI(n22389), .I0(n610_c), .I1(VCC_net), 
            .CO(n22390));
    SB_DFF i890_891 (.Q(n1229), .C(clock_c), .D(n11817));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_195_i1_3_lut (.I0(ootx_payloads_0_80), .I1(ootx_payloads_1_80), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[80]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_195_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_196_i1_3_lut (.I0(ootx_payloads_0_79), .I1(ootx_payloads_1_79), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[79]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_196_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_197_i1_3_lut (.I0(ootx_payloads_0_78), .I1(ootx_payloads_1_78), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[78]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_197_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1674_7_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n22634), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_16 (.CI(n22715), .I0(n2699), .I1(n2720), 
            .CO(n22716));
    SB_LUT4 EnabledDecoder_2_i161_2_lut_3_lut (.I0(n66_adj_1904), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n161));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i161_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_CARRY mod_155_add_2009_6 (.CI(n22758), .I0(n2909), .I1(n25182), 
            .CO(n22759));
    SB_DFF i887_888 (.Q(n1230), .C(clock_c), .D(n11816));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_198_i1_3_lut (.I0(ootx_payloads_0_77), .I1(ootx_payloads_1_77), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[77]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_198_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_370 (.I0(n134_adj_1948), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n838));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_370.LUT_INIT = 16'h0020;
    SB_LUT4 i1_3_lut_adj_371 (.I0(n432), .I1(n1087), .I2(data_counters_N_1776), 
            .I3(GND_net), .O(n24028));
    defparam i1_3_lut_adj_371.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_155_add_1205_16_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n22510), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_7 (.CI(n22634), .I0(n2408), .I1(n2423), 
            .CO(n22635));
    SB_LUT4 mod_155_add_468_4_lut (.I0(GND_net), .I1(n611), .I2(VCC_net), 
            .I3(n22388), .O(n89[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_468_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_from_nskip_rise_640_add_4_5_lut (.I0(n6362), .I1(n2280), 
            .I2(counter_from_nskip_rise[3]), .I3(n22353), .O(n91[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 Mux_199_i1_3_lut (.I0(ootx_payloads_0_76), .I1(ootx_payloads_1_76), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[76]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_199_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i884_885 (.Q(n1231), .C(clock_c), .D(n11815));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1205_16 (.CI(n22510), .I0(n1699), .I1(n1730), 
            .CO(n22511));
    SB_LUT4 mod_155_add_1875_15_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n22714), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7002_3_lut_4_lut (.I0(n704), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_91), .O(n11112));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7002_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_468_4 (.CI(n22388), .I0(n611), .I1(VCC_net), 
            .CO(n22389));
    SB_CARRY counter_from_nskip_rise_640_add_4_5 (.CI(n22353), .I0(n2280), 
            .I1(counter_from_nskip_rise[3]), .CO(n22354));
    SB_LUT4 Mux_200_i1_3_lut (.I0(ootx_payloads_0_75), .I1(ootx_payloads_1_75), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[75]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_200_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i881_882 (.Q(n1232), .C(clock_c), .D(n11814));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7594_3_lut_4_lut (.I0(n704), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1342), .O(n11704));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7594_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7515_3_lut_4_lut (.I0(n546), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1421), .O(n11625));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7515_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2143_21 (.CI(n22830), .I0(n3095), .I1(n3116), 
            .CO(n22831));
    SB_LUT4 i6892_3_lut_4_lut (.I0(n546), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_12), .O(n11002));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6892_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2076_12 (.CI(n22792), .I0(n3003), .I1(n3017), 
            .CO(n22793));
    SB_LUT4 mod_155_add_1674_6_lut (.I0(n2409), .I1(n2409), .I2(n25194), 
            .I3(n22633), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_2143_20_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n22829), .O(n37_adj_1966)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i878_879 (.Q(n1233), .C(clock_c), .D(n11813));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_372 (.I0(n128), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n960));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_372.LUT_INIT = 16'h0080;
    SB_CARRY mod_155_add_2143_20 (.CI(n22829), .I0(n3096), .I1(n3116), 
            .CO(n22830));
    SB_LUT4 mod_155_add_2009_5_lut (.I0(n2910), .I1(n2910), .I2(n2918), 
            .I3(n22757), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 counter_from_nskip_rise_640_add_4_4_lut (.I0(n6363), .I1(n2280), 
            .I2(counter_from_nskip_rise[2]), .I3(n22352), .O(n91[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 Mux_201_i1_3_lut (.I0(ootx_payloads_0_74), .I1(ootx_payloads_1_74), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[74]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_201_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7660_3_lut_4_lut (.I0(n836), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1276), .O(n11770));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7660_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_202_i1_3_lut (.I0(ootx_payloads_0_73), .I1(ootx_payloads_1_73), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[73]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_202_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7068_3_lut_4_lut (.I0(n836), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_157), .O(n11178));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7068_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_203_i1_3_lut (.I0(ootx_payloads_0_72), .I1(ootx_payloads_1_72), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[72]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_203_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i875_876 (.Q(n1234), .C(clock_c), .D(n11812));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7514_3_lut_4_lut (.I0(n544), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1422), .O(n11624));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7514_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1875_15 (.CI(n22714), .I0(n2700), .I1(n2720), 
            .CO(n22715));
    SB_LUT4 i6893_3_lut_4_lut (.I0(n544), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_11), .O(n11003));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_373 (.I0(n132), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n836));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_373.LUT_INIT = 16'h0020;
    SB_CARRY mod_155_add_1674_6 (.CI(n22633), .I0(n2409), .I1(n25194), 
            .CO(n22634));
    SB_CARRY counter_from_nskip_rise_640_add_4_4 (.CI(n22352), .I0(n2280), 
            .I1(counter_from_nskip_rise[2]), .CO(n22353));
    SB_LUT4 mod_155_add_2143_19_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n22828), .O(n35_adj_1958)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i872_873 (.Q(n1235), .C(clock_c), .D(n11811));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7513_3_lut_4_lut (.I0(n542), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1423), .O(n11623));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7513_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6894_3_lut_4_lut (.I0(n542), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_10), .O(n11004));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7659_3_lut_4_lut (.I0(n834), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1277), .O(n11769));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7659_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_15_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n22509), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2143_19 (.CI(n22828), .I0(n3097), .I1(n3116), 
            .CO(n22829));
    SB_LUT4 Mux_204_i1_3_lut (.I0(ootx_payloads_0_71), .I1(ootx_payloads_1_71), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[71]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_204_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7067_3_lut_4_lut (.I0(n834), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_156), .O(n11177));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7067_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_205_i1_3_lut (.I0(ootx_payloads_0_70), .I1(ootx_payloads_1_70), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[70]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_205_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7512_3_lut_4_lut (.I0(n540), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1424), .O(n11622));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7512_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_468_3_lut (.I0(GND_net), .I1(n612_c), .I2(VCC_net), 
            .I3(n22387), .O(n89[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_468_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF i869_870 (.Q(n1236), .C(clock_c), .D(n11810));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i6895_3_lut_4_lut (.I0(n540), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_9), .O(n11005));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6895_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7028_3_lut_4_lut (.I0(n756), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_117), .O(n11138));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7028_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1205_15 (.CI(n22509), .I0(n1700), .I1(n1730), 
            .CO(n22510));
    SB_CARRY mod_155_add_2009_5 (.CI(n22757), .I0(n2910), .I1(n2918), 
            .CO(n22758));
    SB_LUT4 Mux_206_i1_3_lut (.I0(ootx_payloads_0_69), .I1(ootx_payloads_1_69), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[69]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_206_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_34_i1_3_lut_adj_374 (.I0(data_counters_0_4), .I1(data_counters_1_4), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[4] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_34_i1_3_lut_adj_374.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_468_3 (.CI(n22387), .I0(n612_c), .I1(VCC_net), 
            .CO(n22388));
    SB_LUT4 mod_155_add_1875_14_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n22713), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2143_18_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n22827), .O(n33_adj_1956)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_207_i1_3_lut (.I0(ootx_payloads_0_68), .I1(ootx_payloads_1_68), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[68]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_207_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i866_867 (.Q(n1237), .C(clock_c), .D(n11809));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_4_lut (.I0(\ootx_payloads_N_1699[6] ), .I1(\ootx_payloads_N_1699[8] ), 
            .I2(n130_adj_2047), .I3(\ootx_payloads_N_1699[7] ), .O(n578));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 mod_155_add_1674_5_lut (.I0(n2410), .I1(n2410), .I2(n2423), 
            .I3(n22632), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1674_5 (.CI(n22632), .I0(n2410), .I1(n2423), 
            .CO(n22633));
    SB_LUT4 i1_2_lut_4_lut_adj_375 (.I0(\ootx_payloads_N_1699[6] ), .I1(\ootx_payloads_N_1699[8] ), 
            .I2(n130_adj_2047), .I3(\ootx_payloads_N_1699[7] ), .O(n834));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_4_lut_adj_375.LUT_INIT = 16'h1000;
    SB_LUT4 Mux_208_i1_3_lut (.I0(ootx_payloads_0_67), .I1(ootx_payloads_1_67), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[67]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_208_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_209_i1_3_lut (.I0(ootx_payloads_0_66), .I1(ootx_payloads_1_66), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[66]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_209_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_210_i1_3_lut (.I0(ootx_payloads_0_65), .I1(ootx_payloads_1_65), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[65]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_210_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i65_2_lut_3_lut (.I0(n17_adj_1864), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n65_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i65_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mod_155_add_1205_14_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n22508), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 counter_from_nskip_rise_640_add_4_3_lut (.I0(n6364), .I1(n2280), 
            .I2(counter_from_nskip_rise[1]), .I3(n22351), .O(n91[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mod_155_add_2143_18 (.CI(n22827), .I0(n3098), .I1(n3116), 
            .CO(n22828));
    SB_DFF i863_864 (.Q(n1238), .C(clock_c), .D(n11808));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_211_i1_3_lut (.I0(ootx_payloads_0_64), .I1(ootx_payloads_1_64), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[64]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_211_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i66_2_lut_3_lut (.I0(n17_adj_1864), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n66_adj_1904));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i66_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mod_155_add_468_2_lut (.I0(GND_net), .I1(n2851[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n89[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_468_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 lighthouse_counter_639_add_4_2_lut (.I0(GND_net), .I1(new_data), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n129[0])) /* synthesis syn_instantiated=1 */ ;
    defparam lighthouse_counter_639_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7001_3_lut_4_lut (.I0(n702), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_90), .O(n11111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7593_3_lut_4_lut (.I0(n702), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1343), .O(n11703));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7593_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i860_861 (.Q(n1239), .C(clock_c), .D(n11807));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7511_3_lut_4_lut (.I0(n538), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1425), .O(n11621));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7511_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6896_3_lut_4_lut (.I0(n538), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_8), .O(n11006));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6896_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_212_i1_3_lut (.I0(ootx_payloads_0_63), .I1(ootx_payloads_1_63), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[63]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_212_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1205_14 (.CI(n22508), .I0(n1701), .I1(n1730), 
            .CO(n22509));
    SB_CARRY counter_from_nskip_rise_640_add_4_3 (.CI(n22351), .I0(n2280), 
            .I1(counter_from_nskip_rise[1]), .CO(n22352));
    SB_LUT4 i7658_3_lut_4_lut (.I0(n832), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1278), .O(n11768));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7658_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_468_2 (.CI(VCC_net), .I0(n2851[26]), .I1(GND_net), 
            .CO(n22387));
    SB_LUT4 Mux_213_i1_3_lut (.I0(ootx_payloads_0_62), .I1(ootx_payloads_1_62), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[62]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_213_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i857_858 (.Q(n1240), .C(clock_c), .D(n11806));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7066_3_lut_4_lut (.I0(n832), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_155), .O(n11176));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7066_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_214_i1_3_lut (.I0(ootx_payloads_0_61), .I1(ootx_payloads_1_61), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[61]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_214_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7510_3_lut_4_lut (.I0(n536), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1426), .O(n11620));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7510_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1875_14 (.CI(n22713), .I0(n2701), .I1(n2720), 
            .CO(n22714));
    SB_LUT4 mod_155_add_1674_4_lut (.I0(n2411), .I1(n2411), .I2(n2423), 
            .I3(n22631), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7620_3_lut_4_lut (.I0(n756), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1316), .O(n11730));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7620_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_215_i1_3_lut (.I0(ootx_payloads_0_60), .I1(ootx_payloads_1_60), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[60]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_215_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6898_3_lut_4_lut (.I0(n536), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_7), .O(n11008));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6898_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_33_i1_3_lut_adj_376 (.I0(data_counters_0_5), .I1(data_counters_1_5), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[5] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_33_i1_3_lut_adj_376.LUT_INIT = 16'hcaca;
    SB_DFF i854_855 (.Q(n1241), .C(clock_c), .D(n11805));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7010_3_lut_4_lut (.I0(n720), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_99), .O(n11120));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7010_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_377 (.I0(n126_adj_1853), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n958));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_377.LUT_INIT = 16'h0080;
    SB_CARRY mod_155_add_1674_4 (.CI(n22631), .I0(n2411), .I1(n2423), 
            .CO(n22632));
    SB_LUT4 i7602_3_lut_4_lut (.I0(n720), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1334), .O(n11712));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_13_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n22507), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 counter_from_nskip_rise_640_add_4_2_lut (.I0(n6365), .I1(n2280), 
            .I2(counter_from_nskip_rise[0]), .I3(VCC_net), .O(n91[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 Mux_216_i1_3_lut (.I0(ootx_payloads_0_59), .I1(ootx_payloads_1_59), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[59]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_216_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i851_852 (.Q(n1242), .C(clock_c), .D(n11804));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 sensor_state_switch_counter_641_add_4_7_lut (.I0(GND_net), .I1(n2276), 
            .I2(sensor_state_switch_counter[5]), .I3(n22386), .O(n100[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sensor_state_switch_counter_641_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_637_16_lut (.I0(GND_net), .I1(n577[15]), .I2(GND_net), 
            .I3(n22319), .O(n4485[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Mux_217_i1_3_lut (.I0(ootx_payloads_0_58), .I1(ootx_payloads_1_58), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[58]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_217_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1205_13 (.CI(n22507), .I0(n1702), .I1(n1730), 
            .CO(n22508));
    SB_CARRY counter_from_nskip_rise_640_add_4_2 (.CI(VCC_net), .I0(n2280), 
            .I1(counter_from_nskip_rise[0]), .CO(n22351));
    SB_LUT4 Mux_218_i1_3_lut (.I0(ootx_payloads_0_57), .I1(ootx_payloads_1_57), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[57]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_218_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i848_849 (.Q(n1243), .C(clock_c), .D(n11803));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_378 (.I0(n128), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n832));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_378.LUT_INIT = 16'h0020;
    SB_LUT4 sensor_state_switch_counter_641_add_4_6_lut (.I0(GND_net), .I1(n2276), 
            .I2(sensor_state_switch_counter[4]), .I3(n22385), .O(n100[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sensor_state_switch_counter_641_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_637_16 (.CI(n22319), .I0(n577[15]), .I1(GND_net), .CO(n4501));
    SB_LUT4 mod_155_add_1674_3_lut (.I0(n2412), .I1(n2412), .I2(n2423), 
            .I3(n22630), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1875_13_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n22712), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7117_3_lut_4_lut (.I0(n934), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_206), .O(n11227));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7117_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7509_3_lut_4_lut (.I0(n534), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1427), .O(n11619));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7509_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_12_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n22506), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i845_846 (.Q(n1244), .C(clock_c), .D(n11802));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1674_3 (.CI(n22630), .I0(n2412), .I1(n2423), 
            .CO(n22631));
    SB_LUT4 Mux_219_i1_3_lut (.I0(ootx_payloads_0_56), .I1(ootx_payloads_1_56), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[56]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_219_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sensor_state_switch_counter_641_add_4_6 (.CI(n22385), .I0(n2276), 
            .I1(sensor_state_switch_counter[4]), .CO(n22386));
    SB_LUT4 i6900_3_lut_4_lut (.I0(n534), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_6), .O(n11010));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6900_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7657_3_lut_4_lut (.I0(n830), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1279), .O(n11767));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7657_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7574_3_lut_4_lut (.I0(n664), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1362), .O(n11684));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_220_i1_3_lut (.I0(ootx_payloads_0_55), .I1(ootx_payloads_1_55), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[55]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_220_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i842_843 (.Q(n1245), .C(clock_c), .D(n11801));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1205_12 (.CI(n22506), .I0(n1703), .I1(n1730), 
            .CO(n22507));
    SB_LUT4 add_637_15_lut (.I0(GND_net), .I1(n577[14]), .I2(GND_net), 
            .I3(n22318), .O(n4485[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sensor_state_switch_counter_641_add_4_5_lut (.I0(GND_net), .I1(n2276), 
            .I2(sensor_state_switch_counter[3]), .I3(n22384), .O(n100[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sensor_state_switch_counter_641_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7065_3_lut_4_lut (.I0(n830), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_154), .O(n11175));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7065_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_221_i1_3_lut (.I0(ootx_payloads_0_54), .I1(ootx_payloads_1_54), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[54]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_221_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7000_3_lut_4_lut (.I0(n700), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_89), .O(n11110));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7000_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_222_i1_3_lut (.I0(ootx_payloads_0_53), .I1(ootx_payloads_1_53), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[53]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_222_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_2009_4_lut (.I0(n2911), .I1(n2911), .I2(n2918), 
            .I3(n22756), .O(n3010)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_637_15 (.CI(n22318), .I0(n577[14]), .I1(GND_net), .CO(n22319));
    SB_LUT4 i7592_3_lut_4_lut (.I0(n700), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1344), .O(n11702));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7592_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i839_840 (.Q(n1246), .C(clock_c), .D(n11800));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1875_13 (.CI(n22712), .I0(n2702), .I1(n2720), 
            .CO(n22713));
    SB_LUT4 mod_155_add_1674_2_lut (.I0(n2851[8]), .I1(n2851[8]), .I2(n25194), 
            .I3(VCC_net), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_379 (.I0(n126_adj_1853), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n830));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_379.LUT_INIT = 16'h0020;
    SB_LUT4 i7508_3_lut_4_lut (.I0(n532), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1428), .O(n11618));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7508_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_223_i1_3_lut (.I0(ootx_payloads_0_52), .I1(ootx_payloads_1_52), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[52]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_223_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6904_3_lut_4_lut (.I0(n532), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_5), .O(n11014));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6904_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7656_3_lut_4_lut (.I0(n828), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1280), .O(n11766));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7656_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i836_837 (.Q(n1247), .C(clock_c), .D(n11799));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1674_2 (.CI(VCC_net), .I0(n2851[8]), .I1(n25194), 
            .CO(n22630));
    SB_LUT4 i7064_3_lut_4_lut (.I0(n828), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_153), .O(n11174));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7064_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7507_3_lut_4_lut (.I0(n530), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1429), .O(n11617));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7507_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6905_3_lut_4_lut (.I0(n530), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_4), .O(n11015));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6905_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_380 (.I0(n124), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n956));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_380.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_1205_11_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n22505), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_14_lut (.I0(GND_net), .I1(n577[13]), .I2(GND_net), 
            .I3(n22317), .O(n4485[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6999_3_lut_4_lut (.I0(n698), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_88), .O(n11109));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6999_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY sensor_state_switch_counter_641_add_4_5 (.CI(n22384), .I0(n2276), 
            .I1(sensor_state_switch_counter[3]), .CO(n22385));
    SB_DFF i833_834 (.Q(n1248), .C(clock_c), .D(n11798));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7591_3_lut_4_lut (.I0(n698), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1345), .O(n11701));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7591_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_224_i1_3_lut (.I0(ootx_payloads_0_51), .I1(ootx_payloads_1_51), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[51]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_224_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_225_i1_3_lut (.I0(ootx_payloads_0_50), .I1(ootx_payloads_1_50), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[50]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_225_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1205_11 (.CI(n22505), .I0(n1704), .I1(n1730), 
            .CO(n22506));
    SB_CARRY add_637_14 (.CI(n22317), .I0(n577[13]), .I1(GND_net), .CO(n22318));
    SB_LUT4 Mux_226_i1_3_lut (.I0(ootx_payloads_0_49), .I1(ootx_payloads_1_49), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[49]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_226_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i122_2_lut (.I0(n57_adj_2045), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_2046));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i122_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_381 (.I0(n124), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n828));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_381.LUT_INIT = 16'h0020;
    SB_DFF i830_831 (.Q(n1249), .C(clock_c), .D(n11797));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_382 (.I0(n122_adj_2046), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n954));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_382.LUT_INIT = 16'h0080;
    SB_LUT4 i7655_3_lut_4_lut (.I0(n826), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1281), .O(n11765));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7655_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_227_i1_3_lut (.I0(ootx_payloads_0_48), .I1(ootx_payloads_1_48), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[48]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_227_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7063_3_lut_4_lut (.I0(n826), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_152), .O(n11173));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7063_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7506_3_lut_4_lut (.I0(n528), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1430), .O(n11616));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7506_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 sensor_state_switch_counter_641_add_4_4_lut (.I0(GND_net), .I1(n2276), 
            .I2(sensor_state_switch_counter[2]), .I3(n22383), .O(n100[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sensor_state_switch_counter_641_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Mux_228_i1_3_lut (.I0(ootx_payloads_0_47), .I1(ootx_payloads_1_47), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[47]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_228_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1607_24_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n22629), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2076_11_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n22791), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2009_4 (.CI(n22756), .I0(n2911), .I1(n2918), 
            .CO(n22757));
    SB_LUT4 i6982_3_lut_4_lut (.I0(n664), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_71), .O(n11092));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6908_3_lut_4_lut (.I0(n528), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_3), .O(n11018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6908_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_10_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n22504), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7505_3_lut_4_lut (.I0(n526), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1431), .O(n11615));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7505_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY sensor_state_switch_counter_641_add_4_4 (.CI(n22383), .I0(n2276), 
            .I1(sensor_state_switch_counter[2]), .CO(n22384));
    SB_LUT4 mod_155_add_1875_12_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n22711), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6911_3_lut_4_lut (.I0(n526), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_2), .O(n11021));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6911_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_229_i1_3_lut (.I0(ootx_payloads_0_46), .I1(ootx_payloads_1_46), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[46]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_229_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_383 (.I0(n122_adj_2046), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n826));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_383.LUT_INIT = 16'h0020;
    SB_LUT4 i6998_3_lut_4_lut (.I0(n696), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_87), .O(n11108));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1205_10 (.CI(n22504), .I0(n1705), .I1(n1730), 
            .CO(n22505));
    SB_LUT4 mod_155_add_1607_23_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n22628), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_230_i1_3_lut (.I0(ootx_payloads_0_45), .I1(ootx_payloads_1_45), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[45]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_230_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sensor_state_switch_counter_641_add_4_3_lut (.I0(GND_net), .I1(n2276), 
            .I2(sensor_state_switch_counter[1]), .I3(n22382), .O(n100[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sensor_state_switch_counter_641_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7590_3_lut_4_lut (.I0(n696), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1346), .O(n11700));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7590_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7654_3_lut_4_lut (.I0(n824), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1282), .O(n11764));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7654_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_231_i1_3_lut (.I0(ootx_payloads_0_44), .I1(ootx_payloads_1_44), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[44]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_231_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7062_3_lut_4_lut (.I0(n824), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_151), .O(n11172));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7062_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_384 (.I0(n120), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n952));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_384.LUT_INIT = 16'h0080;
    SB_LUT4 Mux_232_i1_3_lut (.I0(ootx_payloads_0_43), .I1(ootx_payloads_1_43), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[43]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_232_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1875_12 (.CI(n22711), .I0(n2703), .I1(n2720), 
            .CO(n22712));
    SB_LUT4 EnabledDecoder_2_i124_2_lut (.I0(n59_adj_1950), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n124));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i124_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7504_3_lut_4_lut (.I0(n524), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1432), .O(n11614));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7504_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1607_23 (.CI(n22628), .I0(n2292), .I1(n2324), 
            .CO(n22629));
    SB_LUT4 add_637_13_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[12] ), 
            .I2(GND_net), .I3(n22316), .O(n4485[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1205_9_lut (.I0(n1706_adj_1810), .I1(n1706_adj_1810), 
            .I2(n1730), .I3(n22503), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6949_3_lut_4_lut (.I0(n524), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_1), .O(n11059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6949_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_233_i1_3_lut (.I0(ootx_payloads_0_42), .I1(ootx_payloads_1_42), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[42]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_233_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_385 (.I0(n120), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n824));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_385.LUT_INIT = 16'h0020;
    SB_LUT4 Mux_234_i1_3_lut (.I0(ootx_payloads_0_41), .I1(ootx_payloads_1_41), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[41]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_234_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sensor_state_switch_counter_641_add_4_3 (.CI(n22382), .I0(n2276), 
            .I1(sensor_state_switch_counter[1]), .CO(n22383));
    SB_CARRY add_637_13 (.CI(n22316), .I0(\ootx_payloads_N_1730[12] ), .I1(GND_net), 
            .CO(n22317));
    SB_LUT4 Mux_235_i1_3_lut (.I0(ootx_payloads_0_40), .I1(ootx_payloads_1_40), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[40]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_235_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_236_i1_3_lut (.I0(ootx_payloads_0_39), .I1(ootx_payloads_1_39), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[39]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_236_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_237_i1_3_lut (.I0(ootx_payloads_0_38), .I1(ootx_payloads_1_38), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[38]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_237_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1205_9 (.CI(n22503), .I0(n1706_adj_1810), .I1(n1730), 
            .CO(n22504));
    SB_LUT4 mod_155_add_1607_22_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n22627), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2143_17_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n22826), .O(n31_adj_1972)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_238_i1_3_lut (.I0(ootx_payloads_0_37), .I1(ootx_payloads_1_37), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[37]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_238_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7503_3_lut_4_lut (.I0(n522), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1433), .O(n11613));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7503_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6950_3_lut_4_lut (.I0(n522), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_0), .O(n11060));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6950_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7653_3_lut_4_lut (.I0(n822), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1283), .O(n11763));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7653_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7061_3_lut_4_lut (.I0(n822), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_150), .O(n11171));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7061_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 sensor_state_switch_counter_641_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(sensor_state_switch_counter[0]), .I3(VCC_net), .O(n100[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sensor_state_switch_counter_641_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6997_3_lut_4_lut (.I0(n694), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_86), .O(n11107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6997_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1607_22 (.CI(n22627), .I0(n2293), .I1(n2324), 
            .CO(n22628));
    SB_LUT4 i7589_3_lut_4_lut (.I0(n694), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1347), .O(n11699));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7589_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_386 (.I0(n118_adj_2055), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n950));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_386.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_1205_8_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n22502), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_12_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[11] ), 
            .I2(GND_net), .I3(n22315), .O(n4485[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sensor_state_switch_counter_641_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(sensor_state_switch_counter[0]), .CO(n22382));
    SB_LUT4 Mux_239_i1_3_lut (.I0(ootx_payloads_0_36), .I1(ootx_payloads_1_36), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[36]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_239_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7018_3_lut_4_lut (.I0(n736), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_107), .O(n11128));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7018_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_240_i1_3_lut (.I0(ootx_payloads_0_35), .I1(ootx_payloads_1_35), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[35]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_240_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7610_3_lut_4_lut (.I0(n736), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1326), .O(n11720));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7610_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6996_3_lut_4_lut (.I0(n692), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_85), .O(n11106));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6996_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1205_8 (.CI(n22502), .I0(n1707), .I1(n1730), 
            .CO(n22503));
    SB_LUT4 Mux_241_i1_3_lut (.I0(ootx_payloads_0_34), .I1(ootx_payloads_1_34), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[34]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_241_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_242_i1_3_lut (.I0(ootx_payloads_0_33), .I1(ootx_payloads_1_33), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[33]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_242_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7588_3_lut_4_lut (.I0(n692), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1348), .O(n11698));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7588_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 counter_from_nskip_rise_640_add_4_33_lut (.I0(n6334), .I1(n2280), 
            .I2(counter_from_nskip_rise[31]), .I3(n22381), .O(n91[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_33_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_637_12 (.CI(n22315), .I0(\ootx_payloads_N_1730[11] ), .I1(GND_net), 
            .CO(n22316));
    SB_LUT4 Mux_243_i1_3_lut (.I0(ootx_payloads_0_32), .I1(ootx_payloads_1_32), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[32]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_243_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_244_i1_3_lut (.I0(ootx_payloads_0_31), .I1(ootx_payloads_1_31), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[31]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_244_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2076_11 (.CI(n22791), .I0(n3004), .I1(n3017), 
            .CO(n22792));
    SB_LUT4 EnabledDecoder_2_i51_2_lut_3_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n51));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i51_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_2009_3_lut (.I0(n2912), .I1(n2912), .I2(n2918), 
            .I3(n22755), .O(n3011)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1875_11_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n22710), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1875_11 (.CI(n22710), .I0(n2704), .I1(n2720), 
            .CO(n22711));
    SB_LUT4 mod_155_add_1607_21_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n22626), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i52_2_lut_3_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n52));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i52_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 Mux_245_i1_3_lut (.I0(ootx_payloads_0_30), .I1(ootx_payloads_1_30), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[30]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_245_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut (.I0(crc32s_N_1751), .I1(ootx_payloads_N_1699[0]), 
            .I2(ootx_payloads_N_1699[1]), .I3(GND_net), .O(n12_adj_2072));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i12_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut (.I0(crc32s_N_1751), .I1(ootx_payloads_N_1699[0]), 
            .I2(ootx_payloads_N_1699[1]), .I3(GND_net), .O(n11_adj_2070));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i11_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY mod_155_add_1607_21 (.CI(n22626), .I0(n2294), .I1(n2324), 
            .CO(n22627));
    SB_CARRY mod_155_add_2143_17 (.CI(n22826), .I0(n3099), .I1(n3116), 
            .CO(n22827));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_387 (.I0(n116), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n948));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_387.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_1205_7_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n22501), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_11_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[10] ), 
            .I2(GND_net), .I3(n22314), .O(n4485[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Mux_246_i1_3_lut (.I0(ootx_payloads_0_29), .I1(ootx_payloads_1_29), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[29]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_246_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_388 (.I0(n118_adj_2055), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n822));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_388.LUT_INIT = 16'h0020;
    SB_LUT4 Mux_247_i1_3_lut (.I0(ootx_payloads_0_28), .I1(ootx_payloads_1_28), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[28]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_247_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_389 (.I0(n2679), .I1(n2680), .I2(n20105), .I3(n3), 
            .O(n1087));
    defparam i3_4_lut_adj_389.LUT_INIT = 16'h0020;
    SB_LUT4 counter_from_nskip_rise_640_add_4_32_lut (.I0(n6335), .I1(n2280), 
            .I2(counter_from_nskip_rise[30]), .I3(n22380), .O(n91[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_32_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mod_155_add_1205_7 (.CI(n22501), .I0(n1708), .I1(n1730), 
            .CO(n22502));
    SB_LUT4 i6995_3_lut_4_lut (.I0(n690), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_84), .O(n11105));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_32 (.CI(n22380), .I0(n2280), 
            .I1(counter_from_nskip_rise[30]), .CO(n22381));
    SB_LUT4 i3_3_lut_adj_390 (.I0(ootx_payloads_N_1744[1]), .I1(n20112), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n22972));
    defparam i3_3_lut_adj_390.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7587_3_lut_4_lut (.I0(n690), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1349), .O(n11697));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7587_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_248_i1_3_lut (.I0(ootx_payloads_0_27), .I1(ootx_payloads_1_27), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[27]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_248_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7027_3_lut_4_lut (.I0(n754), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_116), .O(n11137));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7027_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1607_20_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n22625), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7619_3_lut_4_lut (.I0(n754), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1317), .O(n11729));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_6_lut (.I0(n1709), .I1(n1709), .I2(n25197), 
            .I3(n22500), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_637_11 (.CI(n22314), .I0(\ootx_payloads_N_1730[10] ), .I1(GND_net), 
            .CO(n22315));
    SB_CARRY mod_155_add_1607_20 (.CI(n22625), .I0(n2295), .I1(n2324), 
            .CO(n22626));
    SB_LUT4 i7708_3_lut_4_lut (.I0(n932), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1228), .O(n11818));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7708_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_249_i1_3_lut (.I0(ootx_payloads_0_26), .I1(ootx_payloads_1_26), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[26]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_249_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_from_nskip_rise_640_add_4_31_lut (.I0(n6336), .I1(n2280), 
            .I2(counter_from_nskip_rise[29]), .I3(n22379), .O(n91[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_31_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_391 (.I0(n114_adj_2044), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n946));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_391.LUT_INIT = 16'h0080;
    SB_CARRY mod_155_add_1205_6 (.CI(n22500), .I0(n1709), .I1(n25197), 
            .CO(n22501));
    SB_LUT4 Mux_250_i1_3_lut (.I0(ootx_payloads_0_25), .I1(ootx_payloads_1_25), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[25]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_250_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_251_i1_3_lut (.I0(ootx_payloads_0_24), .I1(ootx_payloads_1_24), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[24]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_251_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_252_i1_3_lut (.I0(ootx_payloads_0_23), .I1(ootx_payloads_1_23), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[23]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_252_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_3_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(GND_net), .O(n63_adj_2059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i63_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut_4_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n96));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i96_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_CARRY counter_from_nskip_rise_640_add_4_31 (.CI(n22379), .I0(n2280), 
            .I1(counter_from_nskip_rise[29]), .CO(n22380));
    SB_LUT4 add_637_10_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[9] ), 
            .I2(GND_net), .I3(n22313), .O(n4485[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut_4_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n95));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i95_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i7573_3_lut_4_lut (.I0(n662), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1363), .O(n11683));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_253_i1_3_lut (.I0(ootx_payloads_0_22), .I1(ootx_payloads_1_22), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[22]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_253_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1875_10_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n22709), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_3_lut_adj_392 (.I0(data_counters_N_1776), .I1(n1087), .I2(n1119), 
            .I3(GND_net), .O(n8_adj_2075));
    defparam i3_3_lut_adj_392.LUT_INIT = 16'hfefe;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n49));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i49_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i50_2_lut_3_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n50));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i50_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i2_2_lut_adj_393 (.I0(ootx_payloads_N_1744[0]), .I1(n20105), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_2077));
    defparam i2_2_lut_adj_393.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_394 (.I0(\lighthouse[0] ), .I1(n9_adj_2077), .I2(n8_adj_2075), 
            .I3(n432), .O(n9771));
    defparam i1_4_lut_adj_394.LUT_INIT = 16'h5554;
    SB_LUT4 i7652_3_lut_4_lut (.I0(n820), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1284), .O(n11762));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7652_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1607_19_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n22624), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_254_i1_3_lut (.I0(ootx_payloads_0_21), .I1(ootx_payloads_1_21), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[21]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_254_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1205_5_lut (.I0(n1710), .I1(n1710), .I2(n1730), 
            .I3(n22499), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 counter_from_nskip_rise_640_add_4_30_lut (.I0(n6337), .I1(n2280), 
            .I2(counter_from_nskip_rise[28]), .I3(n22378), .O(n91[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_30_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_637_10 (.CI(n22313), .I0(\ootx_payloads_N_1730[9] ), .I1(GND_net), 
            .CO(n22314));
    SB_CARRY mod_155_add_1205_5 (.CI(n22499), .I0(n1710), .I1(n1730), 
            .CO(n22500));
    SB_LUT4 i7060_3_lut_4_lut (.I0(n820), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_149), .O(n11170));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7060_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_255_i1_3_lut (.I0(ootx_payloads_0_20), .I1(ootx_payloads_1_20), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[20]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_255_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2009_3 (.CI(n22755), .I0(n2912), .I1(n2918), 
            .CO(n22756));
    SB_LUT4 EnabledDecoder_2_i128_2_lut (.I0(n63_adj_2059), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n128));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i128_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6994_3_lut_4_lut (.I0(n688), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_83), .O(n11104));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6994_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7586_3_lut_4_lut (.I0(n688), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1350), .O(n11696));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7586_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_30 (.CI(n22378), .I0(n2280), 
            .I1(counter_from_nskip_rise[28]), .CO(n22379));
    SB_CARRY mod_155_add_1875_10 (.CI(n22709), .I0(n2705), .I1(n2720), 
            .CO(n22710));
    SB_LUT4 EnabledDecoder_2_i10_2_lut_3_lut (.I0(crc32s_N_1751), .I1(ootx_payloads_N_1699[0]), 
            .I2(ootx_payloads_N_1699[1]), .I3(GND_net), .O(n10_adj_2079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i10_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut (.I0(crc32s_N_1751), .I1(ootx_payloads_N_1699[0]), 
            .I2(ootx_payloads_N_1699[1]), .I3(GND_net), .O(n9));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i9_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_CARRY mod_155_add_1607_19 (.CI(n22624), .I0(n2296), .I1(n2324), 
            .CO(n22625));
    SB_LUT4 mod_155_add_1607_18_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n22623), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_256_i1_3_lut (.I0(ootx_payloads_0_19), .I1(ootx_payloads_1_19), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[19]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_256_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6981_3_lut_4_lut (.I0(n662), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_70), .O(n11091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_257_i1_3_lut (.I0(ootx_payloads_0_18), .I1(ootx_payloads_1_18), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[18]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_257_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_395 (.I0(n116), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n820));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_395.LUT_INIT = 16'h0020;
    SB_LUT4 Mux_258_i1_3_lut (.I0(ootx_payloads_0_17), .I1(ootx_payloads_1_17), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[17]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_258_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1205_4_lut (.I0(n1711), .I1(n1711), .I2(n1730), 
            .I3(n22498), .O(n1810)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_396 (.I0(n112_adj_2043), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n944));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_396.LUT_INIT = 16'h0080;
    SB_LUT4 counter_from_nskip_rise_640_add_4_29_lut (.I0(n6338), .I1(n2280), 
            .I2(counter_from_nskip_rise[27]), .I3(n22377), .O(n91[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_29_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i6993_3_lut_4_lut (.I0(n686), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_82), .O(n11103));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6993_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_259_i1_3_lut (.I0(ootx_payloads_0_16), .I1(ootx_payloads_1_16), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[16]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_259_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7585_3_lut_4_lut (.I0(n686), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1351), .O(n11695));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7585_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1205_4 (.CI(n22498), .I0(n1711), .I1(n1730), 
            .CO(n22499));
    SB_CARRY counter_from_nskip_rise_640_add_4_29 (.CI(n22377), .I0(n2280), 
            .I1(counter_from_nskip_rise[27]), .CO(n22378));
    SB_LUT4 add_637_9_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[8] ), 
            .I2(GND_net), .I3(n22312), .O(n4485[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n47));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i47_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_2009_2_lut (.I0(n2851[3]), .I1(n2851[3]), .I2(n25182), 
            .I3(VCC_net), .O(n3012)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_1875_9_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n22708), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i48_2_lut_3_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n48));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i48_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_CARRY add_637_9 (.CI(n22312), .I0(\ootx_payloads_N_1730[8] ), .I1(GND_net), 
            .CO(n22313));
    SB_LUT4 i7651_3_lut_4_lut (.I0(n818), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1285), .O(n11761));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7651_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_260_i1_3_lut (.I0(ootx_payloads_0_15), .I1(ootx_payloads_1_15), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[15]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_260_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_261_i1_3_lut (.I0(ootx_payloads_0_14), .I1(ootx_payloads_1_14), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[14]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_261_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1607_18 (.CI(n22623), .I0(n2297), .I1(n2324), 
            .CO(n22624));
    SB_LUT4 i7059_3_lut_4_lut (.I0(n818), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_148), .O(n11169));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7059_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_262_i1_3_lut (.I0(ootx_payloads_0_13), .I1(ootx_payloads_1_13), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[13]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_262_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_263_i1_3_lut (.I0(ootx_payloads_0_12), .I1(ootx_payloads_1_12), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[12]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_263_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7116_3_lut_4_lut (.I0(n932), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_205), .O(n11226));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7116_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_3_lut (.I0(n1712), .I1(n1712), .I2(n1730), 
            .I3(n22497), .O(n1811)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_397 (.I0(n110_adj_1911), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n942));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_397.LUT_INIT = 16'h0080;
    SB_LUT4 mod_155_add_1607_17_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n22622), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 counter_from_nskip_rise_640_add_4_28_lut (.I0(n6339), .I1(n2280), 
            .I2(counter_from_nskip_rise[26]), .I3(n22376), .O(n91[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_28_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_398 (.I0(n114_adj_2044), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n818));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_398.LUT_INIT = 16'h0020;
    SB_LUT4 Mux_264_i1_3_lut (.I0(ootx_payloads_0_11), .I1(ootx_payloads_1_11), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[11]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_264_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_1205_3 (.CI(n22497), .I0(n1712), .I1(n1730), 
            .CO(n22498));
    SB_LUT4 EnabledDecoder_2_i130_2_lut (.I0(n65_c), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n130_adj_2047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i130_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY counter_from_nskip_rise_640_add_4_28 (.CI(n22376), .I0(n2280), 
            .I1(counter_from_nskip_rise[26]), .CO(n22377));
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n45));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i45_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i46_2_lut_3_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n46));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i46_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_CARRY mod_155_add_1607_17 (.CI(n22622), .I0(n2298), .I1(n2324), 
            .CO(n22623));
    SB_LUT4 Mux_265_i1_3_lut (.I0(ootx_payloads_0_10), .I1(ootx_payloads_1_10), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[10]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_265_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_637_8_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[7] ), 
            .I2(GND_net), .I3(n22311), .O(n4485[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_399 (.I0(n95), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n992));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_399.LUT_INIT = 16'h0080;
    SB_LUT4 i7650_3_lut_4_lut (.I0(n816), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1286), .O(n11760));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7650_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_266_i1_3_lut (.I0(ootx_payloads_0_9), .I1(ootx_payloads_1_9), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[9]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_266_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7058_3_lut_4_lut (.I0(n816), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_147), .O(n11168));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7058_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1205_2_lut (.I0(n2851[15]), .I1(n2851[15]), .I2(n25197), 
            .I3(VCC_net), .O(n1812)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 counter_from_nskip_rise_640_add_4_27_lut (.I0(n6340), .I1(n2280), 
            .I2(counter_from_nskip_rise[25]), .I3(n22375), .O(n91[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_27_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_637_8 (.CI(n22311), .I0(\ootx_payloads_N_1730[7] ), .I1(GND_net), 
            .CO(n22312));
    SB_LUT4 Mux_267_i1_3_lut (.I0(ootx_payloads_0_8), .I1(ootx_payloads_1_8), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[8]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_267_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7822_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_25), 
            .I3(\ootx_crc32_o[1] [25]), .O(n11932));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7822_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY mod_155_add_1205_2 (.CI(VCC_net), .I0(n2851[15]), .I1(n25197), 
            .CO(n22497));
    SB_LUT4 i7827_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_30), 
            .I3(\ootx_crc32_o[1] [30]), .O(n11937));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7827_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY mod_155_add_1875_9 (.CI(n22708), .I0(n2706), .I1(n2720), 
            .CO(n22709));
    SB_LUT4 i7824_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_27), 
            .I3(\ootx_crc32_o[1] [27]), .O(n11934));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7824_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7823_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_26), 
            .I3(\ootx_crc32_o[1] [26]), .O(n11933));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7823_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7828_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_31), 
            .I3(\ootx_crc32_o[1] [31]), .O(n11938));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7828_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY counter_from_nskip_rise_640_add_4_27 (.CI(n22375), .I0(n2280), 
            .I1(counter_from_nskip_rise[25]), .CO(n22376));
    SB_LUT4 i7826_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_29), 
            .I3(\ootx_crc32_o[1] [29]), .O(n11936));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7826_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7825_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_28), 
            .I3(\ootx_crc32_o[1] [28]), .O(n11935));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7825_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7821_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_24), 
            .I3(\ootx_crc32_o[1] [24]), .O(n11931));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7821_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_1607_16_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n22621), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1875_8_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n22707), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7820_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_23), 
            .I3(\ootx_crc32_o[1] [23]), .O(n11930));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7820_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7819_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_22), 
            .I3(\ootx_crc32_o[1] [22]), .O(n11929));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7819_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7818_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_21), 
            .I3(\ootx_crc32_o[1] [21]), .O(n11928));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7818_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY mod_155_add_1607_16 (.CI(n22621), .I0(n2299), .I1(n2324), 
            .CO(n22622));
    SB_LUT4 Mux_268_i1_3_lut (.I0(ootx_payloads_0_7), .I1(ootx_payloads_1_7), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[7]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_268_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7817_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_20), 
            .I3(\ootx_crc32_o[1] [20]), .O(n11927));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7817_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_1138_17_lut (.I0(n1598_adj_2086), .I1(n1598_adj_2086), 
            .I2(n1631_adj_2058), .I3(n22496), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_7_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[6] ), 
            .I2(GND_net), .I3(n22310), .O(n4485[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7572_3_lut_4_lut (.I0(n660), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1364), .O(n11682));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_269_i1_3_lut (.I0(ootx_payloads_0_6), .I1(ootx_payloads_1_6), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[6]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_269_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_270_i1_3_lut (.I0(ootx_payloads_0_5), .I1(ootx_payloads_1_5), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[5]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_270_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7816_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_19), 
            .I3(\ootx_crc32_o[1] [19]), .O(n11926));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7816_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7815_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_18), 
            .I3(\ootx_crc32_o[1] [18]), .O(n11925));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7815_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7814_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_17), 
            .I3(\ootx_crc32_o[1] [17]), .O(n11924));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7814_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7813_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_16), 
            .I3(\ootx_crc32_o[1] [16]), .O(n11923));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7813_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7812_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_15), 
            .I3(\ootx_crc32_o[1] [15]), .O(n11922));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7812_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 counter_from_nskip_rise_640_add_4_26_lut (.I0(n6341), .I1(n2280), 
            .I2(counter_from_nskip_rise[24]), .I3(n22374), .O(n91[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_26_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i7811_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_14), 
            .I3(\ootx_crc32_o[1] [14]), .O(n11921));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7811_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7810_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_13), 
            .I3(\ootx_crc32_o[1] [13]), .O(n11920));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7810_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_1138_16_lut (.I0(n1599_adj_2087), .I1(n1599_adj_2087), 
            .I2(n1631_adj_2058), .I3(n22495), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_637_7 (.CI(n22310), .I0(\ootx_payloads_N_1730[6] ), .I1(GND_net), 
            .CO(n22311));
    SB_LUT4 i7809_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_12), 
            .I3(\ootx_crc32_o[1] [12]), .O(n11919));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7809_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7808_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_11), 
            .I3(\ootx_crc32_o[1] [11]), .O(n11918));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7808_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7807_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_10), 
            .I3(\ootx_crc32_o[1] [10]), .O(n11917));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7807_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY counter_from_nskip_rise_640_add_4_26 (.CI(n22374), .I0(n2280), 
            .I1(counter_from_nskip_rise[24]), .CO(n22375));
    SB_LUT4 mod_155_add_1607_15_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n22620), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_32_i1_3_lut_adj_400 (.I0(data_counters_0_6), .I1(data_counters_1_6), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[6] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_32_i1_3_lut_adj_400.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_31_i1_3_lut_adj_401 (.I0(data_counters_0_7), .I1(data_counters_1_7), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[7] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_31_i1_3_lut_adj_401.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_30_i1_3_lut_adj_402 (.I0(data_counters_0_8), .I1(data_counters_1_8), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[8] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_30_i1_3_lut_adj_402.LUT_INIT = 16'hcaca;
    SB_LUT4 i7806_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_9), 
            .I3(\ootx_crc32_o[1] [9]), .O(n11916));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7806_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7805_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_8), 
            .I3(\ootx_crc32_o[1] [8]), .O(n11915));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7805_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7804_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_7), 
            .I3(\ootx_crc32_o[1] [7]), .O(n11914));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7804_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7803_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_6), 
            .I3(\ootx_crc32_o[1] [6]), .O(n11913));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7803_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7802_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_5), 
            .I3(\ootx_crc32_o[1] [5]), .O(n11912));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7802_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7801_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_4), 
            .I3(\ootx_crc32_o[1] [4]), .O(n11911));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7801_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7800_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_3), 
            .I3(\ootx_crc32_o[1] [3]), .O(n11910));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7800_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7799_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_2), 
            .I3(\ootx_crc32_o[1] [2]), .O(n11909));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7799_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 Mux_271_i1_3_lut (.I0(ootx_payloads_0_4), .I1(ootx_payloads_1_4), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[4]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_271_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_272_i1_3_lut (.I0(ootx_payloads_0_3), .I1(ootx_payloads_1_3), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[3]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_272_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6902_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_0), 
            .I3(\ootx_crc32_o[1] [0]), .O(n11012));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i6902_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_2143_16_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n22825), .O(n29_adj_1957)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1607_15 (.CI(n22620), .I0(n2300), .I1(n2324), 
            .CO(n22621));
    SB_LUT4 Mux_273_i1_3_lut (.I0(ootx_payloads_0_2), .I1(ootx_payloads_1_2), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[2]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_273_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7798_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(crc32s_1_1), 
            .I3(\ootx_crc32_o[1] [1]), .O(n11908));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7798_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY mod_155_add_2143_16 (.CI(n22825), .I0(n3100), .I1(n3116), 
            .CO(n22826));
    SB_CARRY mod_155_add_1138_16 (.CI(n22495), .I0(n1599_adj_2087), .I1(n1631_adj_2058), 
            .CO(n22496));
    SB_LUT4 add_637_6_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[5] ), 
            .I2(GND_net), .I3(n22309), .O(n4485[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_155_add_2009_2 (.CI(VCC_net), .I0(n2851[3]), .I1(n25182), 
            .CO(n22755));
    SB_LUT4 Mux_274_i1_3_lut (.I0(ootx_payloads_0_1), .I1(ootx_payloads_1_1), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_274_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_2143_15_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n22824), .O(n27_adj_1954)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2076_10_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n22790), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i43_2_lut_3_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n43));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i43_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 Mux_25_i1_3_lut_adj_403 (.I0(bit_counters_0_11), .I1(bit_counters_1_11), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[11]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_25_i1_3_lut_adj_403.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_12_i1_3_lut_adj_404 (.I0(bit_counters_0_24), .I1(bit_counters_1_24), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[24]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_12_i1_3_lut_adj_404.LUT_INIT = 16'hcaca;
    SB_CARRY mod_155_add_2143_15 (.CI(n22824), .I0(n3101), .I1(n3116), 
            .CO(n22825));
    SB_LUT4 counter_from_nskip_rise_640_add_4_25_lut (.I0(n6342), .I1(n2280), 
            .I2(counter_from_nskip_rise[23]), .I3(n22373), .O(n91[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i20512_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25180));
    defparam i20512_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i44_2_lut_3_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n44));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i44_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_405 (.I0(n112_adj_2043), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n816));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_405.LUT_INIT = 16'h0020;
    SB_LUT4 mod_155_add_1138_15_lut (.I0(n1600_adj_2090), .I1(n1600_adj_2090), 
            .I2(n1631_adj_2058), .I3(n22494), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_637_6 (.CI(n22309), .I0(\ootx_payloads_N_1730[5] ), .I1(GND_net), 
            .CO(n22310));
    SB_LUT4 Mux_11_i1_3_lut_adj_406 (.I0(bit_counters_0_25), .I1(bit_counters_1_25), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[25]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_11_i1_3_lut_adj_406.LUT_INIT = 16'hcaca;
    SB_DFF i827_828 (.Q(n1250), .C(clock_c), .D(n11796));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i824_825 (.Q(n1251), .C(clock_c), .D(n11795));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i821_822 (.Q(n1252), .C(clock_c), .D(n11794));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i818_819 (.Q(n1253), .C(clock_c), .D(n11793));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i815_816 (.Q(n1254), .C(clock_c), .D(n11792));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i812_813 (.Q(n1255), .C(clock_c), .D(n11791));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i809_810 (.Q(n1256), .C(clock_c), .D(n11790));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i806_807 (.Q(n1257), .C(clock_c), .D(n11789));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i803_804 (.Q(n1258), .C(clock_c), .D(n11788));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i800_801 (.Q(n1259), .C(clock_c), .D(n11787));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i797_798 (.Q(n1260), .C(clock_c), .D(n11786));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i794_795 (.Q(n1261), .C(clock_c), .D(n11785));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i791_792 (.Q(n1262), .C(clock_c), .D(n11784));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i788_789 (.Q(n1263), .C(clock_c), .D(n11783));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i785_786 (.Q(n1264), .C(clock_c), .D(n11782));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i782_783 (.Q(n1265), .C(clock_c), .D(n11781));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i779_780 (.Q(n1266), .C(clock_c), .D(n11780));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i776_777 (.Q(n1267), .C(clock_c), .D(n11779));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i773_774 (.Q(n1268), .C(clock_c), .D(n11778));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i770_771 (.Q(n1269), .C(clock_c), .D(n11777));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i767_768 (.Q(n1270), .C(clock_c), .D(n11776));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i764_765 (.Q(n1271), .C(clock_c), .D(n11775));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i761_762 (.Q(n1272), .C(clock_c), .D(n11774));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i758_759 (.Q(n1273), .C(clock_c), .D(n11773));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i755_756 (.Q(n1274), .C(clock_c), .D(n11772));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i752_753 (.Q(n1275), .C(clock_c), .D(n11771));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i749_750 (.Q(n1276), .C(clock_c), .D(n11770));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i746_747 (.Q(n1277), .C(clock_c), .D(n11769));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i743_744 (.Q(n1278), .C(clock_c), .D(n11768));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i740_741 (.Q(n1279), .C(clock_c), .D(n11767));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i737_738 (.Q(n1280), .C(clock_c), .D(n11766));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1607_14_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n22619), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_2143_14_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n22823), .O(n25_adj_1953)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i52_3_lut_4_lut (.I0(n13), .I1(n24018), .I2(ootx_payloads_N_1744[1]), 
            .I3(n23974), .O(n22_adj_1846));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i52_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i51_3_lut_4_lut_3_lut (.I0(n13), .I1(n24018), .I2(data), .I3(GND_net), 
            .O(n28));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i51_3_lut_4_lut_3_lut.LUT_INIT = 16'h4e4e;
    SB_LUT4 i1_2_lut_adj_407 (.I0(n2887), .I1(n2900), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_2092));
    defparam i1_2_lut_adj_407.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_408 (.I0(n2897), .I1(n2907), .I2(n2898), .I3(n2889), 
            .O(n42_adj_2093));
    defparam i17_4_lut_adj_408.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_409 (.I0(n2892), .I1(n2893), .I2(n2890), .I3(n2885), 
            .O(n40_adj_2094));
    defparam i15_4_lut_adj_409.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_410 (.I0(n2906), .I1(n2905), .I2(n2896), .I3(n2894), 
            .O(n41_adj_2095));
    defparam i16_4_lut_adj_410.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_411 (.I0(n2908), .I1(n2888), .I2(n2886), .I3(n2901), 
            .O(n39_adj_2096));
    defparam i14_4_lut_adj_411.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_412 (.I0(n2851[3]), .I1(n2912), .I2(n2911), .I3(n2910), 
            .O(n22891));
    defparam i3_4_lut_adj_412.LUT_INIT = 16'hfffe;
    SB_LUT4 i7649_3_lut_4_lut (.I0(n814), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1287), .O(n11759));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7649_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7057_3_lut_4_lut (.I0(n814), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_146), .O(n11167));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7057_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i41_2_lut_3_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n41));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i41_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i42_2_lut_3_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n42));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i42_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_413 (.I0(n110_adj_1911), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n814));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_413.LUT_INIT = 16'h0020;
    SB_LUT4 i6980_3_lut_4_lut (.I0(n660), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_69), .O(n11090));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6980_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i734_735 (.Q(n1281), .C(clock_c), .D(n11765));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i731_732 (.Q(n1282), .C(clock_c), .D(n11764));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i728_729 (.Q(n1283), .C(clock_c), .D(n11763));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i725_726 (.Q(n1284), .C(clock_c), .D(n11762));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i722_723 (.Q(n1285), .C(clock_c), .D(n11761));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i719_720 (.Q(n1286), .C(clock_c), .D(n11760));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i716_717 (.Q(n1287), .C(clock_c), .D(n11759));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i713_714 (.Q(n1288), .C(clock_c), .D(n11758));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i710_711 (.Q(n1289), .C(clock_c), .D(n11757));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i707_708 (.Q(n1290), .C(clock_c), .D(n11756));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i704_705 (.Q(n1291), .C(clock_c), .D(n11755));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i701_702 (.Q(n1292), .C(clock_c), .D(n11754));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i698_699 (.Q(n1293), .C(clock_c), .D(n11753));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i695_696 (.Q(n1294), .C(clock_c), .D(n11752));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i692_693 (.Q(n1295), .C(clock_c), .D(n11751));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i689_690 (.Q(n1296), .C(clock_c), .D(n11750));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i686_687 (.Q(n1297), .C(clock_c), .D(n11749));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i683_684 (.Q(n1298), .C(clock_c), .D(n11748));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i680_681 (.Q(n1299), .C(clock_c), .D(n11747));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i677_678 (.Q(n1300), .C(clock_c), .D(n11746));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i674_675 (.Q(n1301), .C(clock_c), .D(n11745));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i671_672 (.Q(n1302), .C(clock_c), .D(n11744));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i668_669 (.Q(n1303), .C(clock_c), .D(n11743));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i665_666 (.Q(n1304), .C(clock_c), .D(n11742));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i662_663 (.Q(n1305), .C(clock_c), .D(n11741));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i659_660 (.Q(n1306), .C(clock_c), .D(n11740));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i656_657 (.Q(n1307), .C(clock_c), .D(n11739));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i653_654 (.Q(n1308), .C(clock_c), .D(n11738));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i650_651 (.Q(n1309), .C(clock_c), .D(n11737));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i647_648_adj_414 (.Q(n1310), .C(clock_c), .D(n11736));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i644_645_adj_415 (.Q(n1311), .C(clock_c), .D(n11735));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i641_642_adj_416 (.Q(n1312), .C(clock_c), .D(n11734));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i638_639_adj_417 (.Q(n1313), .C(clock_c), .D(n11733));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i635_636_adj_418 (.Q(n1314), .C(clock_c), .D(n11732));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i632_633_adj_419 (.Q(n1315), .C(clock_c), .D(n11731));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i629_630_adj_420 (.Q(n1316), .C(clock_c), .D(n11730));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i626_627_adj_421 (.Q(n1317), .C(clock_c), .D(n11729));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i623_624_adj_422 (.Q(n1318), .C(clock_c), .D(n11728));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i620_621_adj_423 (.Q(n1319), .C(clock_c), .D(n11727));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i617_618_adj_424 (.Q(n1320), .C(clock_c), .D(n11726));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i614_615_adj_425 (.Q(n1321), .C(clock_c), .D(n11725));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i611_612_adj_426 (.Q(n1322), .C(clock_c), .D(n11724));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i608_609_adj_427 (.Q(n1323), .C(clock_c), .D(n11723));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i605_606_adj_428 (.Q(n1324), .C(clock_c), .D(n11722));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i602_603_adj_429 (.Q(n1325), .C(clock_c), .D(n11721));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i599_600_adj_430 (.Q(n1326), .C(clock_c), .D(n11720));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i596_597_adj_431 (.Q(n1327), .C(clock_c), .D(n11719));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i593_594_adj_432 (.Q(n1328), .C(clock_c), .D(n11718));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i590_591_adj_433 (.Q(n1329), .C(clock_c), .D(n11717));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i587_588_adj_434 (.Q(n1330), .C(clock_c), .D(n11716));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i584_585_adj_435 (.Q(n1331), .C(clock_c), .D(n11715));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i581_582_adj_436 (.Q(n1332), .C(clock_c), .D(n11714));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i578_579_adj_437 (.Q(n1333), .C(clock_c), .D(n11713));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i575_576_adj_438 (.Q(n1334), .C(clock_c), .D(n11712));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i572_573_adj_439 (.Q(n1335), .C(clock_c), .D(n11711));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i569_570_adj_440 (.Q(n1336), .C(clock_c), .D(n11710));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i566_567_adj_441 (.Q(n1337), .C(clock_c), .D(n11709));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i563_564_adj_442 (.Q(n1338), .C(clock_c), .D(n11708));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i560_561_adj_443 (.Q(n1339), .C(clock_c), .D(n11707));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i557_558_adj_444 (.Q(n1340), .C(clock_c), .D(n11706));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i554_555_adj_445 (.Q(n1341), .C(clock_c), .D(n11705));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i551_552_adj_446 (.Q(n1342), .C(clock_c), .D(n11704));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i548_549_adj_447 (.Q(n1343), .C(clock_c), .D(n11703));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i545_546_adj_448 (.Q(n1344), .C(clock_c), .D(n11702));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i542_543_adj_449 (.Q(n1345), .C(clock_c), .D(n11701));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i539_540_adj_450 (.Q(n1346), .C(clock_c), .D(n11700));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i536_537_adj_451 (.Q(n1347), .C(clock_c), .D(n11699));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i533_534_adj_452 (.Q(n1348), .C(clock_c), .D(n11698));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i530_531_adj_453 (.Q(n1349), .C(clock_c), .D(n11697));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i527_528_adj_454 (.Q(n1350), .C(clock_c), .D(n11696));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i524_525_adj_455 (.Q(n1351), .C(clock_c), .D(n11695));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i521_522_adj_456 (.Q(n1352), .C(clock_c), .D(n11694));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i518_519_adj_457 (.Q(n1353), .C(clock_c), .D(n11693));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i515_516_adj_458 (.Q(n1354), .C(clock_c), .D(n11692));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i512_513 (.Q(n1355), .C(clock_c), .D(n11691));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i509_510 (.Q(n1356), .C(clock_c), .D(n11690));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i506_507 (.Q(n1357), .C(clock_c), .D(n11689));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i503_504 (.Q(n1358), .C(clock_c), .D(n11688));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i500_501 (.Q(n1359), .C(clock_c), .D(n11687));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i497_498 (.Q(n1360), .C(clock_c), .D(n11686));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i494_495 (.Q(n1361), .C(clock_c), .D(n11685));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i491_492 (.Q(n1362), .C(clock_c), .D(n11684));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i488_489 (.Q(n1363), .C(clock_c), .D(n11683));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i485_486 (.Q(n1364), .C(clock_c), .D(n11682));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i482_483 (.Q(n1365), .C(clock_c), .D(n11681));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i479_480 (.Q(n1366), .C(clock_c), .D(n11680));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i476_477 (.Q(n1367), .C(clock_c), .D(n11679));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i473_474 (.Q(n1368), .C(clock_c), .D(n11678));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i470_471 (.Q(n1369), .C(clock_c), .D(n11677));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i467_468 (.Q(n1370), .C(clock_c), .D(n11676));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i464_465 (.Q(n1371), .C(clock_c), .D(n11675));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i461_462 (.Q(n1372), .C(clock_c), .D(n11674));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i458_459 (.Q(n1373), .C(clock_c), .D(n11673));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i455_456 (.Q(n1374), .C(clock_c), .D(n11672));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i452_453 (.Q(n1375), .C(clock_c), .D(n11671));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i449_450 (.Q(n1376), .C(clock_c), .D(n11670));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i446_447 (.Q(n1377), .C(clock_c), .D(n11669));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i443_444 (.Q(n1378), .C(clock_c), .D(n11668));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i440_441 (.Q(n1379), .C(clock_c), .D(n11667));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i437_438 (.Q(n1380), .C(clock_c), .D(n11666));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i434_435 (.Q(n1381), .C(clock_c), .D(n11665));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i431_432 (.Q(n1382), .C(clock_c), .D(n11664));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i428_429 (.Q(n1383), .C(clock_c), .D(n11663));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i425_426 (.Q(n1384), .C(clock_c), .D(n11662));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i422_423 (.Q(n1385), .C(clock_c), .D(n11661));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i419_420 (.Q(n1386), .C(clock_c), .D(n11660));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i416_417 (.Q(n1387), .C(clock_c), .D(n11659));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i413_414 (.Q(n1388), .C(clock_c), .D(n11658));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i410_411 (.Q(n1389), .C(clock_c), .D(n11657));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i407_408 (.Q(n1390), .C(clock_c), .D(n11656));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i404_405 (.Q(n1391), .C(clock_c), .D(n11655));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i401_402 (.Q(n1392), .C(clock_c), .D(n11654));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i398_399 (.Q(n1393), .C(clock_c), .D(n11653));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i395_396 (.Q(n1394), .C(clock_c), .D(n11652));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i392_393 (.Q(n1395), .C(clock_c), .D(n11651));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i389_390 (.Q(n1396), .C(clock_c), .D(n11650));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i386_387 (.Q(n1397), .C(clock_c), .D(n11649));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i383_384 (.Q(n1398), .C(clock_c), .D(n11648));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i380_381 (.Q(n1399), .C(clock_c), .D(n11647));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i377_378 (.Q(n1400), .C(clock_c), .D(n11646));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i374_375 (.Q(n1401), .C(clock_c), .D(n11645));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i371_372 (.Q(n1402), .C(clock_c), .D(n11644));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i368_369 (.Q(n1403), .C(clock_c), .D(n11643));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i365_366 (.Q(n1404), .C(clock_c), .D(n11642));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i362_363 (.Q(n1405), .C(clock_c), .D(n11641));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i359_360 (.Q(n1406), .C(clock_c), .D(n11640));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i356_357 (.Q(n1407), .C(clock_c), .D(n11639));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i353_354 (.Q(n1408), .C(clock_c), .D(n11638));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i350_351 (.Q(n1409), .C(clock_c), .D(n11637));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i347_348 (.Q(n1410), .C(clock_c), .D(n11636));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i344_345 (.Q(n1411), .C(clock_c), .D(n11635));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i341_342 (.Q(n1412), .C(clock_c), .D(n11634));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i338_339 (.Q(n1413), .C(clock_c), .D(n11633));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i335_336 (.Q(n1414), .C(clock_c), .D(n11632));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i332_333 (.Q(n1415), .C(clock_c), .D(n11631));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i329_330 (.Q(n1416), .C(clock_c), .D(n11630));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i326_327 (.Q(n1417), .C(clock_c), .D(n11629));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i323_324 (.Q(n1418), .C(clock_c), .D(n11628));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i320_321 (.Q(n1419), .C(clock_c), .D(n11627));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i317_318 (.Q(n1420), .C(clock_c), .D(n11626));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i314_315 (.Q(n1421), .C(clock_c), .D(n11625));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i311_312 (.Q(n1422), .C(clock_c), .D(n11624));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i308_309 (.Q(n1423), .C(clock_c), .D(n11623));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i305_306 (.Q(n1424), .C(clock_c), .D(n11622));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i302_303 (.Q(n1425), .C(clock_c), .D(n11621));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i299_300 (.Q(n1426), .C(clock_c), .D(n11620));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i296_297 (.Q(n1427), .C(clock_c), .D(n11619));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i293_294 (.Q(n1428), .C(clock_c), .D(n11618));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i290_291 (.Q(n1429), .C(clock_c), .D(n11617));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i287_288 (.Q(n1430), .C(clock_c), .D(n11616));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i284_285 (.Q(n1431), .C(clock_c), .D(n11615));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i281_282 (.Q(n1432), .C(clock_c), .D(n11614));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i278_279 (.Q(n1433), .C(clock_c), .D(n11613));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i131_132 (.Q(n3112[31]), .C(clock_c), .D(n11612));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i128_129_adj_459 (.Q(n3112[30]), .C(clock_c), .D(n11611));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i125_126 (.Q(n3112[29]), .C(clock_c), .D(n11610));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i122_123 (.Q(n3112[28]), .C(clock_c), .D(n11609));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i119_120 (.Q(n3112[27]), .C(clock_c), .D(n11608));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i116_117_adj_460 (.Q(n3112[26]), .C(clock_c), .D(n11607));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i113_114 (.Q(n3112[25]), .C(clock_c), .D(n11606));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i110_111 (.Q(n3112[24]), .C(clock_c), .D(n11605));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i107_108 (.Q(n3112[23]), .C(clock_c), .D(n11604));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i104_105_adj_461 (.Q(n3112[22]), .C(clock_c), .D(n22997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i101_102 (.Q(n3112[21]), .C(clock_c), .D(n11602));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i98_99 (.Q(n3112[20]), .C(clock_c), .D(n23001));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i95_96 (.Q(n3112[19]), .C(clock_c), .D(n11600));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i92_93_adj_462 (.Q(n3112[18]), .C(clock_c), .D(n11599));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i89_90 (.Q(n3112[17]), .C(clock_c), .D(n11598));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i86_87 (.Q(n3112[16]), .C(clock_c), .D(n11597));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i83_84 (.Q(n3112[15]), .C(clock_c), .D(n11596));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i80_81_adj_463 (.Q(n3112[14]), .C(clock_c), .D(n11595));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i77_78 (.Q(n3112[13]), .C(clock_c), .D(n11594));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i74_75 (.Q(n3112[12]), .C(clock_c), .D(n11593));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i71_72 (.Q(n3112[11]), .C(clock_c), .D(n11592));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i68_69_adj_464 (.Q(n3112[10]), .C(clock_c), .D(n11591));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i65_66 (.Q(n3112[9]), .C(clock_c), .D(n11590));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i62_63 (.Q(n3112[8]), .C(clock_c), .D(n11589));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i59_60 (.Q(n3112[7]), .C(clock_c), .D(n11588));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i56_57_adj_465 (.Q(n3112[6]), .C(clock_c), .D(n11587));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i53_54 (.Q(n3112[5]), .C(clock_c), .D(n11586));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i50_51 (.Q(n3112[4]), .C(clock_c), .D(n11585));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i47_48 (.Q(n3112[3]), .C(clock_c), .D(n11584));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i44_45_adj_466 (.Q(n3112[2]), .C(clock_c), .D(n11583));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i41_42 (.Q(n3112[1]), .C(clock_c), .D(n11582));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i38_39 (.Q(n3112[0]), .C(clock_c), .D(n11581));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i227_228 (.Q(crc32s_1_31), .C(clock_c), .D(n11580));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i224_225 (.Q(crc32s_1_30), .C(clock_c), .D(n11579));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i221_222 (.Q(crc32s_1_29), .C(clock_c), .D(n11578));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i218_219 (.Q(crc32s_1_28), .C(clock_c), .D(n11577));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i215_216 (.Q(crc32s_1_27), .C(clock_c), .D(n11576));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i212_213 (.Q(crc32s_1_26), .C(clock_c), .D(n11575));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i209_210 (.Q(crc32s_1_25), .C(clock_c), .D(n11574));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i206_207 (.Q(crc32s_1_24), .C(clock_c), .D(n11573));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i203_204 (.Q(crc32s_1_23), .C(clock_c), .D(n11572));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i200_201 (.Q(crc32s_1_22), .C(clock_c), .D(n11571));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i197_198 (.Q(crc32s_1_21), .C(clock_c), .D(n11570));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i194_195 (.Q(crc32s_1_20), .C(clock_c), .D(n11569));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i191_192 (.Q(crc32s_1_19), .C(clock_c), .D(n11568));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i188_189 (.Q(crc32s_1_18), .C(clock_c), .D(n11567));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i185_186 (.Q(crc32s_1_17), .C(clock_c), .D(n11566));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i182_183 (.Q(crc32s_1_16), .C(clock_c), .D(n11565));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i179_180 (.Q(crc32s_1_15), .C(clock_c), .D(n11564));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i176_177 (.Q(crc32s_1_14), .C(clock_c), .D(n11563));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i173_174 (.Q(crc32s_1_13), .C(clock_c), .D(n11562));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i170_171 (.Q(crc32s_1_12), .C(clock_c), .D(n11561));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i167_168 (.Q(crc32s_1_11), .C(clock_c), .D(n11560));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i164_165 (.Q(crc32s_1_10), .C(clock_c), .D(n11559));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i161_162 (.Q(crc32s_1_9), .C(clock_c), .D(n11558));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i158_159 (.Q(crc32s_1_8), .C(clock_c), .D(n11557));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i155_156 (.Q(crc32s_1_7), .C(clock_c), .D(n11556));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i152_153 (.Q(crc32s_1_6), .C(clock_c), .D(n11555));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i149_150 (.Q(crc32s_1_5), .C(clock_c), .D(n11554));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i146_147 (.Q(crc32s_1_4), .C(clock_c), .D(n11553));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i143_144 (.Q(crc32s_1_3), .C(clock_c), .D(n11552));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i140_141_adj_467 (.Q(crc32s_1_2), .C(clock_c), .D(n11551));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i137_138 (.Q(crc32s_1_1), .C(clock_c), .D(n11550));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i134_135 (.Q(crc32s_1_0), .C(clock_c), .D(n11549));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(49[9:15])
    SB_DFF i1883_1884 (.Q(ootx_payloads_1_263), .C(clock_c), .D(n11548));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1880_1881 (.Q(ootx_payloads_1_262), .C(clock_c), .D(n11547));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1877_1878 (.Q(ootx_payloads_1_261), .C(clock_c), .D(n11546));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1874_1875 (.Q(ootx_payloads_1_260), .C(clock_c), .D(n11545));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1871_1872 (.Q(ootx_payloads_1_259), .C(clock_c), .D(n11544));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1868_1869 (.Q(ootx_payloads_1_258), .C(clock_c), .D(n11543));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1865_1866 (.Q(ootx_payloads_1_257), .C(clock_c), .D(n11542));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1862_1863 (.Q(ootx_payloads_1_256), .C(clock_c), .D(n11541));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1859_1860 (.Q(ootx_payloads_1_255), .C(clock_c), .D(n11540));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1856_1857 (.Q(ootx_payloads_1_254), .C(clock_c), .D(n11539));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1853_1854 (.Q(ootx_payloads_1_253), .C(clock_c), .D(n11538));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1850_1851 (.Q(ootx_payloads_1_252), .C(clock_c), .D(n11537));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1847_1848 (.Q(ootx_payloads_1_251), .C(clock_c), .D(n11536));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1844_1845 (.Q(ootx_payloads_1_250), .C(clock_c), .D(n11535));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1841_1842 (.Q(ootx_payloads_1_249), .C(clock_c), .D(n11534));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1838_1839 (.Q(ootx_payloads_1_248), .C(clock_c), .D(n11533));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1835_1836 (.Q(ootx_payloads_1_247), .C(clock_c), .D(n11532));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1832_1833 (.Q(ootx_payloads_1_246), .C(clock_c), .D(n11531));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1829_1830 (.Q(ootx_payloads_1_245), .C(clock_c), .D(n11530));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1826_1827 (.Q(ootx_payloads_1_244), .C(clock_c), .D(n11529));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1823_1824 (.Q(ootx_payloads_1_243), .C(clock_c), .D(n11528));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1820_1821 (.Q(ootx_payloads_1_242), .C(clock_c), .D(n11527));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1817_1818 (.Q(ootx_payloads_1_241), .C(clock_c), .D(n11526));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1814_1815 (.Q(ootx_payloads_1_240), .C(clock_c), .D(n11525));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1811_1812 (.Q(ootx_payloads_1_239), .C(clock_c), .D(n11524));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1808_1809 (.Q(ootx_payloads_1_238), .C(clock_c), .D(n11523));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1805_1806 (.Q(ootx_payloads_1_237), .C(clock_c), .D(n11522));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1802_1803 (.Q(ootx_payloads_1_236), .C(clock_c), .D(n11521));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1799_1800 (.Q(ootx_payloads_1_235), .C(clock_c), .D(n11520));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1796_1797 (.Q(ootx_payloads_1_234), .C(clock_c), .D(n11519));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1793_1794 (.Q(ootx_payloads_1_233), .C(clock_c), .D(n11518));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1790_1791 (.Q(ootx_payloads_1_232), .C(clock_c), .D(n11517));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1787_1788 (.Q(ootx_payloads_1_231), .C(clock_c), .D(n11516));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1784_1785 (.Q(ootx_payloads_1_230), .C(clock_c), .D(n11515));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1781_1782 (.Q(ootx_payloads_1_229), .C(clock_c), .D(n11514));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1778_1779 (.Q(ootx_payloads_1_228), .C(clock_c), .D(n11513));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1775_1776 (.Q(ootx_payloads_1_227), .C(clock_c), .D(n11512));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1772_1773 (.Q(ootx_payloads_1_226), .C(clock_c), .D(n11511));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1769_1770 (.Q(ootx_payloads_1_225), .C(clock_c), .D(n11510));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1766_1767 (.Q(ootx_payloads_1_224), .C(clock_c), .D(n11509));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1763_1764 (.Q(ootx_payloads_1_223), .C(clock_c), .D(n11508));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1760_1761 (.Q(ootx_payloads_1_222), .C(clock_c), .D(n11507));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1757_1758 (.Q(ootx_payloads_1_221), .C(clock_c), .D(n11506));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1754_1755 (.Q(ootx_payloads_1_220), .C(clock_c), .D(n11505));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1751_1752 (.Q(ootx_payloads_1_219), .C(clock_c), .D(n11504));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n39));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i39_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i7571_3_lut_4_lut (.I0(n658), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1365), .O(n11681));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n40));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i6979_3_lut_4_lut (.I0(n658), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_68), .O(n11089));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7648_3_lut_4_lut (.I0(n812), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1288), .O(n11758));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7648_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7056_3_lut_4_lut (.I0(n812), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_145), .O(n11166));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7056_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_2_lut (.I0(n2904), .I1(n2903), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_2133));
    defparam i11_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7720_3_lut_4_lut (.I0(n956), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1216), .O(n11830));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7720_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_25 (.CI(n22373), .I0(n2280), 
            .I1(counter_from_nskip_rise[23]), .CO(n22374));
    SB_CARRY mod_155_add_2143_14 (.CI(n22823), .I0(n3102), .I1(n3116), 
            .CO(n22824));
    SB_LUT4 EnabledDecoder_2_i37_2_lut_3_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n37));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i37_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[3] ), 
            .O(n38));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i38_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i6930_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_16), .I3(ootx_shift_registers_0_17), 
            .O(n11040));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6930_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2143_13_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n22822), .O(n23_adj_1974)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6925_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_11), .I3(ootx_shift_registers_0_12), 
            .O(n11035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6925_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6920_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_6), .I3(ootx_shift_registers_0_7), 
            .O(n11030));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6920_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6929_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_15), .I3(ootx_shift_registers_0_16), 
            .O(n11039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6929_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2076_10 (.CI(n22790), .I0(n3005), .I1(n3017), 
            .CO(n22791));
    SB_LUT4 mod_155_add_2076_9_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n22789), .O(n3105_adj_2136)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6916_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_2), .I3(ootx_shift_registers_0_3), 
            .O(n11026));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6916_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6924_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_10), .I3(ootx_shift_registers_0_11), 
            .O(n11034));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6924_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1942_29_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n22754), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_28_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n22753), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_24_i1_3_lut_adj_468 (.I0(bit_counters_0_12), .I1(bit_counters_1_12), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[12]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_24_i1_3_lut_adj_468.LUT_INIT = 16'hcaca;
    SB_LUT4 i6921_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_7), .I3(ootx_shift_registers_0_8), 
            .O(n11031));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6921_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6915_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_1), .I3(ootx_shift_registers_0_2), 
            .O(n11025));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6915_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6923_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_9), .I3(ootx_shift_registers_0_10), 
            .O(n11033));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6923_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6922_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_8), .I3(ootx_shift_registers_0_9), 
            .O(n11032));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6922_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6914_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_0), .I3(ootx_shift_registers_0_1), 
            .O(n11024));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6914_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6913_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(data), .I3(ootx_shift_registers_0_0), .O(n11023));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6913_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7128_3_lut_4_lut (.I0(n956), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_217), .O(n11238));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7128_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6927_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_13), .I3(ootx_shift_registers_0_14), 
            .O(n11037));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6927_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6918_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_4), .I3(ootx_shift_registers_0_5), 
            .O(n11028));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6918_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6926_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_12), .I3(ootx_shift_registers_0_13), 
            .O(n11036));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6926_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1875_8 (.CI(n22707), .I0(n2707), .I1(n2720), 
            .CO(n22708));
    SB_LUT4 mod_155_add_1875_7_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n22706), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6919_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_5), .I3(ootx_shift_registers_0_6), 
            .O(n11029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6919_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1607_14 (.CI(n22619), .I0(n2301), .I1(n2324), 
            .CO(n22620));
    SB_LUT4 mod_155_add_1607_13_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n22618), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19_4_lut_adj_469 (.I0(n2895), .I1(n2899), .I2(n2891), .I3(n26_adj_2092), 
            .O(n44_adj_2137));
    defparam i19_4_lut_adj_469.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_470 (.I0(n39_adj_2096), .I1(n41_adj_2095), .I2(n40_adj_2094), 
            .I3(n42_adj_2093), .O(n48_adj_2138));
    defparam i23_4_lut_adj_470.LUT_INIT = 16'hfffe;
    SB_LUT4 i6928_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_14), .I3(ootx_shift_registers_0_15), 
            .O(n11038));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6928_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6917_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_0_3), .I3(ootx_shift_registers_0_4), 
            .O(n11027));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(89[42:45])
    defparam i6917_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7570_3_lut_4_lut (.I0(n656), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1366), .O(n11680));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7796_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[30]), 
            .I3(\ootx_crc32_o[0] [30]), .O(n11906));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7796_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7795_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[29]), 
            .I3(\ootx_crc32_o[0] [29]), .O(n11905));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7795_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7794_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[28]), 
            .I3(\ootx_crc32_o[0] [28]), .O(n11904));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7794_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7789_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[23]), 
            .I3(\ootx_crc32_o[0] [23]), .O(n11899));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7789_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7793_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[27]), 
            .I3(\ootx_crc32_o[0] [27]), .O(n11903));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7793_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7791_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[25]), 
            .I3(\ootx_crc32_o[0] [25]), .O(n11901));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7791_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7790_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[24]), 
            .I3(\ootx_crc32_o[0] [24]), .O(n11900));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7790_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7792_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[26]), 
            .I3(\ootx_crc32_o[0] [26]), .O(n11902));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7792_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7797_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[31]), 
            .I3(\ootx_crc32_o[0] [31]), .O(n11907));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7797_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14679_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[22]), 
            .I3(\ootx_crc32_o[0] [22]), .O(n11898));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i14679_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7787_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[21]), 
            .I3(\ootx_crc32_o[0] [21]), .O(n11897));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7787_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14639_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[20]), 
            .I3(\ootx_crc32_o[0] [20]), .O(n11896));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i14639_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7785_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[19]), 
            .I3(\ootx_crc32_o[0] [19]), .O(n11895));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7785_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6978_3_lut_4_lut (.I0(n656), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_67), .O(n11088));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6978_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7784_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[18]), 
            .I3(\ootx_crc32_o[0] [18]), .O(n11894));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7784_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14598_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[17]), 
            .I3(\ootx_crc32_o[0] [17]), .O(n11893));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i14598_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7782_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[16]), 
            .I3(\ootx_crc32_o[0] [16]), .O(n11892));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7782_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7781_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[15]), 
            .I3(\ootx_crc32_o[0] [15]), .O(n11891));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7781_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7780_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[14]), 
            .I3(\ootx_crc32_o[0] [14]), .O(n11890));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7780_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7779_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[13]), 
            .I3(\ootx_crc32_o[0] [13]), .O(n11889));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7779_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7778_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[12]), 
            .I3(\ootx_crc32_o[0] [12]), .O(n11888));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7778_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY mod_155_add_1138_15 (.CI(n22494), .I0(n1600_adj_2090), .I1(n1631_adj_2058), 
            .CO(n22495));
    SB_LUT4 i7777_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[11]), 
            .I3(\ootx_crc32_o[0] [11]), .O(n11887));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7777_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7776_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[10]), 
            .I3(\ootx_crc32_o[0] [10]), .O(n11886));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7776_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 counter_from_nskip_rise_640_add_4_24_lut (.I0(n6343), .I1(n2280), 
            .I2(counter_from_nskip_rise[22]), .I3(n22372), .O(n91[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i7775_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[9]), 
            .I3(\ootx_crc32_o[0] [9]), .O(n11885));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7775_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7774_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[8]), 
            .I3(\ootx_crc32_o[0] [8]), .O(n11884));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7774_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7719_3_lut_4_lut (.I0(n954), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1217), .O(n11829));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7719_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7773_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[7]), 
            .I3(\ootx_crc32_o[0] [7]), .O(n11883));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7773_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i20511_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25179));
    defparam i20511_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7772_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[6]), 
            .I3(\ootx_crc32_o[0] [6]), .O(n11882));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7772_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_2_lut_adj_471 (.I0(n1405_c), .I1(n1403_c), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_2139));
    defparam i2_2_lut_adj_471.LUT_INIT = 16'heeee;
    SB_LUT4 i7771_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[5]), 
            .I3(\ootx_crc32_o[0] [5]), .O(n11881));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7771_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_472 (.I0(n2851[18]), .I1(n1412_c), .I2(n1411_c), 
            .I3(n1410_c), .O(n22868));
    defparam i3_4_lut_adj_472.LUT_INIT = 16'hfffe;
    SB_LUT4 i7770_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[4]), 
            .I3(\ootx_crc32_o[0] [4]), .O(n11880));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7770_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7769_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[3]), 
            .I3(\ootx_crc32_o[0] [3]), .O(n11879));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7769_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7768_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[2]), 
            .I3(\ootx_crc32_o[0] [2]), .O(n11878));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7768_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6901_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[0]), 
            .I3(\ootx_crc32_o[0] [0]), .O(n11011));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i6901_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7767_3_lut_4_lut (.I0(\lighthouse[0] ), .I1(n20123), .I2(n3112[1]), 
            .I3(\ootx_crc32_o[0] [1]), .O(n11877));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(85[28:46])
    defparam i7767_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7647_3_lut_4_lut (.I0(n810), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1289), .O(n11757));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7647_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7055_3_lut_4_lut (.I0(n810), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_144), .O(n11165));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7055_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7646_3_lut_4_lut (.I0(n808), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1290), .O(n11756));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7054_3_lut_4_lut (.I0(n808), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_143), .O(n11164));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7054_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut (.I0(n19263), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n17));
    defparam EnabledDecoder_2_i36_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i15371_2_lut_3_lut (.I0(n19263), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n19468));
    defparam i15371_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 EnabledDecoder_2_i16_2_lut_3_lut_4_lut (.I0(ootx_payloads_N_1699[0]), 
            .I1(n88), .I2(ootx_payloads_N_1699[2]), .I3(ootx_payloads_N_1699[1]), 
            .O(n16_adj_2143));
    defparam EnabledDecoder_2_i16_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 EnabledDecoder_2_i17_2_lut_3_lut_4_lut_adj_473 (.I0(ootx_payloads_N_1699[0]), 
            .I1(n88), .I2(ootx_payloads_N_1699[2]), .I3(ootx_payloads_N_1699[1]), 
            .O(n17_adj_2144));
    defparam EnabledDecoder_2_i17_2_lut_3_lut_4_lut_adj_473.LUT_INIT = 16'h0100;
    SB_LUT4 i7645_3_lut_4_lut (.I0(n806), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1291), .O(n11755));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7645_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7053_3_lut_4_lut (.I0(n806), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_142), .O(n11163));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7053_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7766_3_lut_4_lut (.I0(n535), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1170), .O(n11876));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7766_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7174_3_lut_4_lut (.I0(n535), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_263), .O(n11284));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7174_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_474 (.I0(n88_adj_1877), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n792));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_474.LUT_INIT = 16'h0020;
    SB_LUT4 i6_4_lut_adj_475 (.I0(n22868), .I1(n12_adj_2139), .I2(n1401_c), 
            .I3(n1409_c), .O(n16_adj_2146));
    defparam i6_4_lut_adj_475.LUT_INIT = 16'hfefc;
    SB_LUT4 i7644_3_lut_4_lut (.I0(n804), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1292), .O(n11754));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7052_3_lut_4_lut (.I0(n804), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_141), .O(n11162));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7052_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_476 (.I0(n1402_c), .I1(n1406_c), .I2(n1407_c), 
            .I3(n1404_c), .O(n17_adj_2147));
    defparam i7_4_lut_adj_476.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_477 (.I0(n17_adj_2147), .I1(n1408_c), .I2(n16_adj_2146), 
            .I3(n1400_c), .O(n1433_c));
    defparam i9_4_lut_adj_477.LUT_INIT = 16'hfffe;
    SB_LUT4 i7765_3_lut_4_lut (.I0(n533), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1171), .O(n11875));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7765_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7173_3_lut_4_lut (.I0(n533), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_262), .O(n11283));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7173_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE counter_from_nskip_rise_640__i1 (.Q(counter_from_nskip_rise[1]), 
            .C(clock_c), .E(n2282), .D(n91[1]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFER led_i0_i1 (.Q(led_c_0), .C(clock_c), .E(n23775), .D(n4731), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i19417_2_lut_4_lut (.I0(n15_adj_2148), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24069));
    defparam i19417_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_LUT4 i19431_2_lut_4_lut (.I0(n15_adj_2148), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24097));
    defparam i19431_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 EnabledDecoder_2_i14_2_lut_3_lut (.I0(n6_adj_2054), .I1(ootx_payloads_N_1699[1]), 
            .I2(ootx_payloads_N_1699[2]), .I3(GND_net), .O(n14_adj_2149));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(119[37:62])
    defparam EnabledDecoder_2_i14_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i15_2_lut_3_lut (.I0(n6_adj_2054), .I1(ootx_payloads_N_1699[1]), 
            .I2(ootx_payloads_N_1699[2]), .I3(GND_net), .O(n15_adj_2148));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(119[37:62])
    defparam EnabledDecoder_2_i15_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_478 (.I0(n86_adj_1860), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n790));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_478.LUT_INIT = 16'h0020;
    SB_DFFER led_i0_i2 (.Q(led_c_1), .C(clock_c), .E(n23995), .D(n9989), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFER led_i0_i3 (.Q(led_c_2), .C(clock_c), .E(n23996), .D(n9989), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFER led_i0_i4 (.Q(led_c_3), .C(clock_c), .E(n23994), .D(n9989), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFER led_i0_i5 (.Q(led_c_4), .C(clock_c), .E(n23991), .D(n9989), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFER led_i0_i6 (.Q(led_c_5), .C(clock_c), .E(n23992), .D(n9989), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFFER led_i0_i7 (.Q(led_c_6), .C(clock_c), .E(n23990), .D(n9989), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF i512_513_adj_479 (.Q(ootx_payloads_0_78), .C(clock_c), .D(n11099));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i509_510_adj_480 (.Q(ootx_payloads_0_77), .C(clock_c), .D(n11098));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7643_3_lut_4_lut (.I0(n802), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1293), .O(n11753));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2076_9 (.CI(n22789), .I0(n3006), .I1(n3017), 
            .CO(n22790));
    SB_LUT4 mod_155_add_1138_14_lut (.I0(n1601_adj_2150), .I1(n1601_adj_2150), 
            .I2(n1631_adj_2058), .I3(n22493), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_5_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[4] ), 
            .I2(GND_net), .I3(n22308), .O(n4485[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7051_3_lut_4_lut (.I0(n802), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_140), .O(n11161));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7051_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_24 (.CI(n22372), .I0(n2280), 
            .I1(counter_from_nskip_rise[22]), .CO(n22373));
    SB_LUT4 i7642_3_lut_4_lut (.I0(n800), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1294), .O(n11752));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7050_3_lut_4_lut (.I0(n800), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_139), .O(n11160));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7050_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19416_2_lut_4_lut (.I0(n17_adj_2144), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24067));
    defparam i19416_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_CARRY mod_155_add_2143_13 (.CI(n22822), .I0(n3103), .I1(n3116), 
            .CO(n22823));
    SB_LUT4 mod_155_add_2143_12_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n22821), .O(n21_adj_1970)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1607_13 (.CI(n22618), .I0(n2302), .I1(n2324), 
            .CO(n22619));
    SB_CARRY add_637_5 (.CI(n22308), .I0(\ootx_payloads_N_1730[4] ), .I1(GND_net), 
            .CO(n22309));
    SB_LUT4 i19457_2_lut_4_lut (.I0(n17_adj_2144), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24124));
    defparam i19457_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 i7764_3_lut_4_lut (.I0(n531), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1172), .O(n11874));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7764_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i506_507_adj_481 (.Q(ootx_payloads_0_76), .C(clock_c), .D(n11097));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i503_504_adj_482 (.Q(ootx_payloads_0_75), .C(clock_c), .D(n11096));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i500_501_adj_483 (.Q(ootx_payloads_0_74), .C(clock_c), .D(n11095));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i497_498_adj_484 (.Q(ootx_payloads_0_73), .C(clock_c), .D(n11094));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i494_495_adj_485 (.Q(ootx_payloads_0_72), .C(clock_c), .D(n11093));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i491_492_adj_486 (.Q(ootx_payloads_0_71), .C(clock_c), .D(n11092));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i488_489_adj_487 (.Q(ootx_payloads_0_70), .C(clock_c), .D(n11091));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i485_486_adj_488 (.Q(ootx_payloads_0_69), .C(clock_c), .D(n11090));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i482_483_adj_489 (.Q(ootx_payloads_0_68), .C(clock_c), .D(n11089));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i479_480_adj_490 (.Q(ootx_payloads_0_67), .C(clock_c), .D(n11088));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i476_477_adj_491 (.Q(ootx_payloads_0_66), .C(clock_c), .D(n11087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i473_474_adj_492 (.Q(ootx_payloads_0_65), .C(clock_c), .D(n11086));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i470_471_adj_493 (.Q(ootx_payloads_0_64), .C(clock_c), .D(n11085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i467_468_adj_494 (.Q(ootx_payloads_0_63), .C(clock_c), .D(n11084));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i464_465_adj_495 (.Q(ootx_payloads_0_62), .C(clock_c), .D(n11083));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i461_462_adj_496 (.Q(ootx_payloads_0_61), .C(clock_c), .D(n11082));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i458_459_adj_497 (.Q(ootx_payloads_0_60), .C(clock_c), .D(n11081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i455_456_adj_498 (.Q(ootx_payloads_0_59), .C(clock_c), .D(n11080));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i452_453_adj_499 (.Q(ootx_payloads_0_58), .C(clock_c), .D(n11079));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i449_450_adj_500 (.Q(ootx_payloads_0_57), .C(clock_c), .D(n11078));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i446_447_adj_501 (.Q(ootx_payloads_0_56), .C(clock_c), .D(n11077));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i443_444_adj_502 (.Q(ootx_payloads_0_55), .C(clock_c), .D(n11076));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i440_441_adj_503 (.Q(ootx_payloads_0_54), .C(clock_c), .D(n11075));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i437_438_adj_504 (.Q(ootx_payloads_0_53), .C(clock_c), .D(n11074));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i434_435_adj_505 (.Q(ootx_payloads_0_52), .C(clock_c), .D(n11073));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i431_432_adj_506 (.Q(ootx_payloads_0_51), .C(clock_c), .D(n11072));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i428_429_adj_507 (.Q(ootx_payloads_0_50), .C(clock_c), .D(n11071));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i425_426_adj_508 (.Q(ootx_payloads_0_49), .C(clock_c), .D(n11070));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i422_423_adj_509 (.Q(ootx_payloads_0_48), .C(clock_c), .D(n11069));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i419_420_adj_510 (.Q(ootx_payloads_0_47), .C(clock_c), .D(n11068));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i416_417_adj_511 (.Q(ootx_payloads_0_46), .C(clock_c), .D(n11067));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i413_414_adj_512 (.Q(ootx_payloads_0_45), .C(clock_c), .D(n11066));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFE counter_from_nskip_rise_640__i2 (.Q(counter_from_nskip_rise[2]), 
            .C(clock_c), .E(n2282), .D(n91[2]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i3 (.Q(counter_from_nskip_rise[3]), 
            .C(clock_c), .E(n2282), .D(n91[3]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i4 (.Q(counter_from_nskip_rise[4]), 
            .C(clock_c), .E(n2282), .D(n91[4]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i5 (.Q(counter_from_nskip_rise[5]), 
            .C(clock_c), .E(n2282), .D(n91[5]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i6 (.Q(counter_from_nskip_rise[6]), 
            .C(clock_c), .E(n2282), .D(n91[6]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i7 (.Q(counter_from_nskip_rise[7]), 
            .C(clock_c), .E(n2282), .D(n91[7]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i8 (.Q(counter_from_nskip_rise[8]), 
            .C(clock_c), .E(n2282), .D(n91[8]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i9 (.Q(counter_from_nskip_rise[9]), 
            .C(clock_c), .E(n2282), .D(n91[9]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i10 (.Q(counter_from_nskip_rise[10]), 
            .C(clock_c), .E(n2282), .D(n91[10]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i11 (.Q(counter_from_nskip_rise[11]), 
            .C(clock_c), .E(n2282), .D(n91[11]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i12 (.Q(counter_from_nskip_rise[12]), 
            .C(clock_c), .E(n2282), .D(n91[12]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i13 (.Q(counter_from_nskip_rise[13]), 
            .C(clock_c), .E(n2282), .D(n91[13]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i14 (.Q(counter_from_nskip_rise[14]), 
            .C(clock_c), .E(n2282), .D(n91[14]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i15 (.Q(counter_from_nskip_rise[15]), 
            .C(clock_c), .E(n2282), .D(n91[15]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i16 (.Q(counter_from_nskip_rise[16]), 
            .C(clock_c), .E(n2282), .D(n91[16]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i17 (.Q(counter_from_nskip_rise[17]), 
            .C(clock_c), .E(n2282), .D(n91[17]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i18 (.Q(counter_from_nskip_rise[18]), 
            .C(clock_c), .E(n2282), .D(n91[18]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i19 (.Q(counter_from_nskip_rise[19]), 
            .C(clock_c), .E(n2282), .D(n91[19]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i20 (.Q(counter_from_nskip_rise[20]), 
            .C(clock_c), .E(n2282), .D(n91[20]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i21 (.Q(counter_from_nskip_rise[21]), 
            .C(clock_c), .E(n2282), .D(n91[21]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i22 (.Q(counter_from_nskip_rise[22]), 
            .C(clock_c), .E(n2282), .D(n91[22]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i23 (.Q(counter_from_nskip_rise[23]), 
            .C(clock_c), .E(n2282), .D(n91[23]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i24 (.Q(counter_from_nskip_rise[24]), 
            .C(clock_c), .E(n2282), .D(n91[24]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i25 (.Q(counter_from_nskip_rise[25]), 
            .C(clock_c), .E(n2282), .D(n91[25]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i26 (.Q(counter_from_nskip_rise[26]), 
            .C(clock_c), .E(n2282), .D(n91[26]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i27 (.Q(counter_from_nskip_rise[27]), 
            .C(clock_c), .E(n2282), .D(n91[27]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i28 (.Q(counter_from_nskip_rise[28]), 
            .C(clock_c), .E(n2282), .D(n91[28]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i29 (.Q(counter_from_nskip_rise[29]), 
            .C(clock_c), .E(n2282), .D(n91[29]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i30 (.Q(counter_from_nskip_rise[30]), 
            .C(clock_c), .E(n2282), .D(n91[30]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFFE counter_from_nskip_rise_640__i31 (.Q(counter_from_nskip_rise[31]), 
            .C(clock_c), .E(n2282), .D(n91[31]));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/vhdl_packages/numeric_std.vhd(1241[12:13])
    SB_DFF i1748_1749 (.Q(ootx_payloads_1_218), .C(clock_c), .D(n11503));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1745_1746 (.Q(ootx_payloads_1_217), .C(clock_c), .D(n11502));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1742_1743 (.Q(ootx_payloads_1_216), .C(clock_c), .D(n11501));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1739_1740 (.Q(ootx_payloads_1_215), .C(clock_c), .D(n11500));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1736_1737 (.Q(ootx_payloads_1_214), .C(clock_c), .D(n11499));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1733_1734 (.Q(ootx_payloads_1_213), .C(clock_c), .D(n11498));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1730_1731 (.Q(ootx_payloads_1_212), .C(clock_c), .D(n11497));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1727_1728 (.Q(ootx_payloads_1_211), .C(clock_c), .D(n11496));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1724_1725 (.Q(ootx_payloads_1_210), .C(clock_c), .D(n11495));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1721_1722 (.Q(ootx_payloads_1_209), .C(clock_c), .D(n11494));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1718_1719 (.Q(ootx_payloads_1_208), .C(clock_c), .D(n11493));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1715_1716 (.Q(ootx_payloads_1_207), .C(clock_c), .D(n11492));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1712_1713 (.Q(ootx_payloads_1_206), .C(clock_c), .D(n11491));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1709_1710 (.Q(ootx_payloads_1_205), .C(clock_c), .D(n11490));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1706_1707 (.Q(ootx_payloads_1_204), .C(clock_c), .D(n11489));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1703_1704 (.Q(ootx_payloads_1_203), .C(clock_c), .D(n11488));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1700_1701 (.Q(ootx_payloads_1_202), .C(clock_c), .D(n11487));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1697_1698 (.Q(ootx_payloads_1_201), .C(clock_c), .D(n11486));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1694_1695 (.Q(ootx_payloads_1_200), .C(clock_c), .D(n11485));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1691_1692 (.Q(ootx_payloads_1_199), .C(clock_c), .D(n11484));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1688_1689 (.Q(ootx_payloads_1_198), .C(clock_c), .D(n11483));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1685_1686 (.Q(ootx_payloads_1_197), .C(clock_c), .D(n11482));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1682_1683 (.Q(ootx_payloads_1_196), .C(clock_c), .D(n11481));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1679_1680 (.Q(ootx_payloads_1_195), .C(clock_c), .D(n11480));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1676_1677 (.Q(ootx_payloads_1_194), .C(clock_c), .D(n11479));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1673_1674 (.Q(ootx_payloads_1_193), .C(clock_c), .D(n11478));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1670_1671 (.Q(ootx_payloads_1_192), .C(clock_c), .D(n11477));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1667_1668 (.Q(ootx_payloads_1_191), .C(clock_c), .D(n11476));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1664_1665 (.Q(ootx_payloads_1_190), .C(clock_c), .D(n11475));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1661_1662 (.Q(ootx_payloads_1_189), .C(clock_c), .D(n11474));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1658_1659 (.Q(ootx_payloads_1_188), .C(clock_c), .D(n11473));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1655_1656 (.Q(ootx_payloads_1_187), .C(clock_c), .D(n11472));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7172_3_lut_4_lut (.I0(n531), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_261), .O(n11282));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7172_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_20_i1_3_lut_adj_513 (.I0(data_counters_0_18), .I1(data_counters_1_18), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1699[18]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_20_i1_3_lut_adj_513.LUT_INIT = 16'hcaca;
    SB_LUT4 ootx_payloads_N_1744_0__bdd_4_lut (.I0(ootx_payloads_N_1744[0]), 
            .I1(n24564), .I2(n28), .I3(ootx_payloads_N_1744[1]), .O(n25219));
    defparam ootx_payloads_N_1744_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_514 (.I0(n84), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n788));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_514.LUT_INIT = 16'h0020;
    SB_DFF i1652_1653 (.Q(ootx_payloads_1_186), .C(clock_c), .D(n11471));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1649_1650 (.Q(ootx_payloads_1_185), .C(clock_c), .D(n11470));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1646_1647 (.Q(ootx_payloads_1_184), .C(clock_c), .D(n11469));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1643_1644 (.Q(ootx_payloads_1_183), .C(clock_c), .D(n11468));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i410_411_adj_515 (.Q(ootx_payloads_0_44), .C(clock_c), .D(n11065));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i407_408_adj_516 (.Q(ootx_payloads_0_43), .C(clock_c), .D(n11064));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i404_405_adj_517 (.Q(ootx_payloads_0_42), .C(clock_c), .D(n11063));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i401_402_adj_518 (.Q(ootx_payloads_0_41), .C(clock_c), .D(n11062));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i398_399_adj_519 (.Q(ootx_payloads_0_40), .C(clock_c), .D(n11061));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1640_1641 (.Q(ootx_payloads_1_182), .C(clock_c), .D(n11467));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1637_1638 (.Q(ootx_payloads_1_181), .C(clock_c), .D(n11466));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1634_1635 (.Q(ootx_payloads_1_180), .C(clock_c), .D(n11465));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1631_1632 (.Q(ootx_payloads_1_179), .C(clock_c), .D(n11464));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1628_1629 (.Q(ootx_payloads_1_178), .C(clock_c), .D(n11463));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1625_1626 (.Q(ootx_payloads_1_177), .C(clock_c), .D(n11462));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1622_1623 (.Q(ootx_payloads_1_176), .C(clock_c), .D(n11461));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1619_1620 (.Q(ootx_payloads_1_175), .C(clock_c), .D(n11460));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1616_1617 (.Q(ootx_payloads_1_174), .C(clock_c), .D(n11459));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1613_1614 (.Q(ootx_payloads_1_173), .C(clock_c), .D(n11458));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1610_1611 (.Q(ootx_payloads_1_172), .C(clock_c), .D(n11457));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1607_1608 (.Q(ootx_payloads_1_171), .C(clock_c), .D(n11456));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1604_1605 (.Q(ootx_payloads_1_170), .C(clock_c), .D(n11455));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1601_1602 (.Q(ootx_payloads_1_169), .C(clock_c), .D(n11454));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1598_1599 (.Q(ootx_payloads_1_168), .C(clock_c), .D(n11453));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1595_1596 (.Q(ootx_payloads_1_167), .C(clock_c), .D(n11452));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1592_1593 (.Q(ootx_payloads_1_166), .C(clock_c), .D(n11451));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1589_1590 (.Q(ootx_payloads_1_165), .C(clock_c), .D(n11450));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1586_1587 (.Q(ootx_payloads_1_164), .C(clock_c), .D(n11449));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1583_1584 (.Q(ootx_payloads_1_163), .C(clock_c), .D(n11448));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1580_1581 (.Q(ootx_payloads_1_162), .C(clock_c), .D(n11447));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1577_1578 (.Q(ootx_payloads_1_161), .C(clock_c), .D(n11446));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1574_1575 (.Q(ootx_payloads_1_160), .C(clock_c), .D(n11445));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1571_1572 (.Q(ootx_payloads_1_159), .C(clock_c), .D(n11444));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1568_1569 (.Q(ootx_payloads_1_158), .C(clock_c), .D(n11443));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1565_1566 (.Q(ootx_payloads_1_157), .C(clock_c), .D(n11442));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1562_1563 (.Q(ootx_payloads_1_156), .C(clock_c), .D(n11441));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1559_1560 (.Q(ootx_payloads_1_155), .C(clock_c), .D(n11440));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1556_1557 (.Q(ootx_payloads_1_154), .C(clock_c), .D(n11439));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1553_1554 (.Q(ootx_payloads_1_153), .C(clock_c), .D(n11438));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1550_1551 (.Q(ootx_payloads_1_152), .C(clock_c), .D(n11437));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1547_1548 (.Q(ootx_payloads_1_151), .C(clock_c), .D(n11436));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1544_1545 (.Q(ootx_payloads_1_150), .C(clock_c), .D(n11435));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1541_1542 (.Q(ootx_payloads_1_149), .C(clock_c), .D(n11434));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1538_1539 (.Q(ootx_payloads_1_148), .C(clock_c), .D(n11433));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1535_1536 (.Q(ootx_payloads_1_147), .C(clock_c), .D(n11432));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1532_1533 (.Q(ootx_payloads_1_146), .C(clock_c), .D(n11431));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1529_1530 (.Q(ootx_payloads_1_145), .C(clock_c), .D(n11430));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1526_1527 (.Q(ootx_payloads_1_144), .C(clock_c), .D(n11429));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1523_1524 (.Q(ootx_payloads_1_143), .C(clock_c), .D(n11428));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1520_1521 (.Q(ootx_payloads_1_142), .C(clock_c), .D(n11427));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1517_1518 (.Q(ootx_payloads_1_141), .C(clock_c), .D(n11426));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1514_1515 (.Q(ootx_payloads_1_140), .C(clock_c), .D(n11425));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1511_1512 (.Q(ootx_payloads_1_139), .C(clock_c), .D(n11424));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1508_1509 (.Q(ootx_payloads_1_138), .C(clock_c), .D(n11423));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1505_1506 (.Q(ootx_payloads_1_137), .C(clock_c), .D(n11422));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1502_1503 (.Q(ootx_payloads_1_136), .C(clock_c), .D(n11421));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1499_1500 (.Q(ootx_payloads_1_135), .C(clock_c), .D(n11420));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1496_1497 (.Q(ootx_payloads_1_134), .C(clock_c), .D(n11419));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1493_1494 (.Q(ootx_payloads_1_133), .C(clock_c), .D(n11418));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1490_1491 (.Q(ootx_payloads_1_132), .C(clock_c), .D(n11417));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1487_1488 (.Q(ootx_payloads_1_131), .C(clock_c), .D(n11416));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1484_1485 (.Q(ootx_payloads_1_130), .C(clock_c), .D(n11415));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1481_1482 (.Q(ootx_payloads_1_129), .C(clock_c), .D(n11414));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1478_1479 (.Q(ootx_payloads_1_128), .C(clock_c), .D(n11413));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1475_1476 (.Q(ootx_payloads_1_127), .C(clock_c), .D(n11412));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1472_1473 (.Q(ootx_payloads_1_126), .C(clock_c), .D(n11411));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1469_1470 (.Q(ootx_payloads_1_125), .C(clock_c), .D(n11410));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1466_1467 (.Q(ootx_payloads_1_124), .C(clock_c), .D(n11409));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1463_1464 (.Q(ootx_payloads_1_123), .C(clock_c), .D(n11408));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1460_1461 (.Q(ootx_payloads_1_122), .C(clock_c), .D(n11407));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1457_1458 (.Q(ootx_payloads_1_121), .C(clock_c), .D(n11406));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1454_1455 (.Q(ootx_payloads_1_120), .C(clock_c), .D(n11405));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1451_1452 (.Q(ootx_payloads_1_119), .C(clock_c), .D(n11404));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1448_1449 (.Q(ootx_payloads_1_118), .C(clock_c), .D(n11403));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1445_1446 (.Q(ootx_payloads_1_117), .C(clock_c), .D(n11402));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1442_1443 (.Q(ootx_payloads_1_116), .C(clock_c), .D(n11401));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1439_1440 (.Q(ootx_payloads_1_115), .C(clock_c), .D(n11400));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1436_1437 (.Q(ootx_payloads_1_114), .C(clock_c), .D(n11399));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1433_1434 (.Q(ootx_payloads_1_113), .C(clock_c), .D(n11398));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1430_1431 (.Q(ootx_payloads_1_112), .C(clock_c), .D(n11397));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1427_1428 (.Q(ootx_payloads_1_111), .C(clock_c), .D(n11396));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1424_1425 (.Q(ootx_payloads_1_110), .C(clock_c), .D(n11395));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1421_1422 (.Q(ootx_payloads_1_109), .C(clock_c), .D(n11394));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1418_1419 (.Q(ootx_payloads_1_108), .C(clock_c), .D(n11393));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1415_1416 (.Q(ootx_payloads_1_107), .C(clock_c), .D(n11392));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1412_1413 (.Q(ootx_payloads_1_106), .C(clock_c), .D(n11391));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1409_1410 (.Q(ootx_payloads_1_105), .C(clock_c), .D(n11390));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1406_1407 (.Q(ootx_payloads_1_104), .C(clock_c), .D(n11389));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1403_1404 (.Q(ootx_payloads_1_103), .C(clock_c), .D(n11388));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1400_1401 (.Q(ootx_payloads_1_102), .C(clock_c), .D(n11387));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1397_1398 (.Q(ootx_payloads_1_101), .C(clock_c), .D(n11386));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1394_1395 (.Q(ootx_payloads_1_100), .C(clock_c), .D(n11385));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1391_1392 (.Q(ootx_payloads_1_99), .C(clock_c), .D(n11384));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1388_1389 (.Q(ootx_payloads_1_98), .C(clock_c), .D(n11383));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1385_1386 (.Q(ootx_payloads_1_97), .C(clock_c), .D(n11382));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1382_1383 (.Q(ootx_payloads_1_96), .C(clock_c), .D(n11381));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1379_1380 (.Q(ootx_payloads_1_95), .C(clock_c), .D(n11380));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1376_1377 (.Q(ootx_payloads_1_94), .C(clock_c), .D(n11379));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1373_1374 (.Q(ootx_payloads_1_93), .C(clock_c), .D(n11378));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1370_1371 (.Q(ootx_payloads_1_92), .C(clock_c), .D(n11377));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1367_1368 (.Q(ootx_payloads_1_91), .C(clock_c), .D(n11376));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1364_1365 (.Q(ootx_payloads_1_90), .C(clock_c), .D(n11375));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1361_1362 (.Q(ootx_payloads_1_89), .C(clock_c), .D(n11374));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1358_1359 (.Q(ootx_payloads_1_88), .C(clock_c), .D(n11373));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1355_1356 (.Q(ootx_payloads_1_87), .C(clock_c), .D(n11372));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1352_1353 (.Q(ootx_payloads_1_86), .C(clock_c), .D(n11371));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1349_1350 (.Q(ootx_payloads_1_85), .C(clock_c), .D(n11370));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1346_1347 (.Q(ootx_payloads_1_84), .C(clock_c), .D(n11369));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1343_1344 (.Q(ootx_payloads_1_83), .C(clock_c), .D(n11368));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1340_1341 (.Q(ootx_payloads_1_82), .C(clock_c), .D(n11367));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1337_1338 (.Q(ootx_payloads_1_81), .C(clock_c), .D(n11366));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1334_1335 (.Q(ootx_payloads_1_80), .C(clock_c), .D(n11365));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1331_1332 (.Q(ootx_payloads_1_79), .C(clock_c), .D(n11364));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1328_1329 (.Q(ootx_payloads_1_78), .C(clock_c), .D(n11363));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1325_1326 (.Q(ootx_payloads_1_77), .C(clock_c), .D(n11362));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1322_1323 (.Q(ootx_payloads_1_76), .C(clock_c), .D(n11361));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1319_1320 (.Q(ootx_payloads_1_75), .C(clock_c), .D(n11360));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1316_1317 (.Q(ootx_payloads_1_74), .C(clock_c), .D(n11359));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1313_1314 (.Q(ootx_payloads_1_73), .C(clock_c), .D(n11358));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1310_1311 (.Q(ootx_payloads_1_72), .C(clock_c), .D(n11357));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1307_1308 (.Q(ootx_payloads_1_71), .C(clock_c), .D(n11356));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1304_1305 (.Q(ootx_payloads_1_70), .C(clock_c), .D(n11355));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1301_1302 (.Q(ootx_payloads_1_69), .C(clock_c), .D(n11354));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1298_1299 (.Q(ootx_payloads_1_68), .C(clock_c), .D(n11353));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1295_1296 (.Q(ootx_payloads_1_67), .C(clock_c), .D(n11352));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1292_1293 (.Q(ootx_payloads_1_66), .C(clock_c), .D(n11351));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1289_1290 (.Q(ootx_payloads_1_65), .C(clock_c), .D(n11350));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1286_1287 (.Q(ootx_payloads_1_64), .C(clock_c), .D(n11349));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1283_1284 (.Q(ootx_payloads_1_63), .C(clock_c), .D(n11348));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1280_1281 (.Q(ootx_payloads_1_62), .C(clock_c), .D(n11347));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1277_1278 (.Q(ootx_payloads_1_61), .C(clock_c), .D(n11346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1274_1275 (.Q(ootx_payloads_1_60), .C(clock_c), .D(n11345));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1271_1272 (.Q(ootx_payloads_1_59), .C(clock_c), .D(n11344));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1268_1269 (.Q(ootx_payloads_1_58), .C(clock_c), .D(n11343));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1265_1266 (.Q(ootx_payloads_1_57), .C(clock_c), .D(n11342));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1262_1263 (.Q(ootx_payloads_1_56), .C(clock_c), .D(n11341));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1259_1260 (.Q(ootx_payloads_1_55), .C(clock_c), .D(n11340));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1256_1257 (.Q(ootx_payloads_1_54), .C(clock_c), .D(n11339));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1253_1254 (.Q(ootx_payloads_1_53), .C(clock_c), .D(n11338));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1250_1251 (.Q(ootx_payloads_1_52), .C(clock_c), .D(n11337));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1247_1248 (.Q(ootx_payloads_1_51), .C(clock_c), .D(n11336));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1244_1245 (.Q(ootx_payloads_1_50), .C(clock_c), .D(n11335));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1241_1242 (.Q(ootx_payloads_1_49), .C(clock_c), .D(n11334));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1238_1239 (.Q(ootx_payloads_1_48), .C(clock_c), .D(n11333));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1235_1236 (.Q(ootx_payloads_1_47), .C(clock_c), .D(n11332));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1232_1233 (.Q(ootx_payloads_1_46), .C(clock_c), .D(n11331));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1229_1230 (.Q(ootx_payloads_1_45), .C(clock_c), .D(n11330));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1226_1227 (.Q(ootx_payloads_1_44), .C(clock_c), .D(n11329));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1223_1224 (.Q(ootx_payloads_1_43), .C(clock_c), .D(n11328));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1220_1221 (.Q(ootx_payloads_1_42), .C(clock_c), .D(n11327));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1217_1218 (.Q(ootx_payloads_1_41), .C(clock_c), .D(n11326));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1214_1215 (.Q(ootx_payloads_1_40), .C(clock_c), .D(n11325));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1211_1212 (.Q(ootx_payloads_1_39), .C(clock_c), .D(n11324));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1208_1209 (.Q(ootx_payloads_1_38), .C(clock_c), .D(n11323));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1205_1206 (.Q(ootx_payloads_1_37), .C(clock_c), .D(n11322));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1202_1203 (.Q(ootx_payloads_1_36), .C(clock_c), .D(n11321));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1199_1200 (.Q(ootx_payloads_1_35), .C(clock_c), .D(n11320));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1196_1197 (.Q(ootx_payloads_1_34), .C(clock_c), .D(n11319));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1193_1194 (.Q(ootx_payloads_1_33), .C(clock_c), .D(n11318));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1190_1191 (.Q(ootx_payloads_1_32), .C(clock_c), .D(n11317));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1187_1188 (.Q(ootx_payloads_1_31), .C(clock_c), .D(n11316));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1184_1185 (.Q(ootx_payloads_1_30), .C(clock_c), .D(n11315));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1181_1182 (.Q(ootx_payloads_1_29), .C(clock_c), .D(n11314));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1178_1179 (.Q(ootx_payloads_1_28), .C(clock_c), .D(n11313));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1175_1176 (.Q(ootx_payloads_1_27), .C(clock_c), .D(n11312));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1172_1173 (.Q(ootx_payloads_1_26), .C(clock_c), .D(n11311));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1169_1170 (.Q(ootx_payloads_1_25), .C(clock_c), .D(n11310));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1166_1167 (.Q(ootx_payloads_1_24), .C(clock_c), .D(n11309));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1163_1164 (.Q(ootx_payloads_1_23), .C(clock_c), .D(n11308));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1160_1161 (.Q(ootx_payloads_1_22), .C(clock_c), .D(n11307));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1157_1158 (.Q(ootx_payloads_1_21), .C(clock_c), .D(n11306));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1154_1155 (.Q(ootx_payloads_1_20), .C(clock_c), .D(n11305));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1151_1152 (.Q(ootx_payloads_1_19), .C(clock_c), .D(n11304));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1148_1149 (.Q(ootx_payloads_1_18), .C(clock_c), .D(n11303));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1145_1146 (.Q(ootx_payloads_1_17), .C(clock_c), .D(n11302));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1142_1143 (.Q(ootx_payloads_1_16), .C(clock_c), .D(n11301));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1139_1140 (.Q(ootx_payloads_1_15), .C(clock_c), .D(n11300));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1136_1137 (.Q(ootx_payloads_1_14), .C(clock_c), .D(n11299));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1133_1134 (.Q(ootx_payloads_1_13), .C(clock_c), .D(n11298));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1130_1131 (.Q(ootx_payloads_1_12), .C(clock_c), .D(n11297));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1127_1128 (.Q(ootx_payloads_1_11), .C(clock_c), .D(n11296));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1124_1125 (.Q(ootx_payloads_1_10), .C(clock_c), .D(n11295));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1121_1122 (.Q(ootx_payloads_1_9), .C(clock_c), .D(n11294));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1118_1119 (.Q(ootx_payloads_1_8), .C(clock_c), .D(n11293));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1115_1116 (.Q(ootx_payloads_1_7), .C(clock_c), .D(n11292));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1112_1113 (.Q(ootx_payloads_1_6), .C(clock_c), .D(n11291));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1109_1110 (.Q(ootx_payloads_1_5), .C(clock_c), .D(n11290));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1106_1107 (.Q(ootx_payloads_1_4), .C(clock_c), .D(n11289));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1103_1104 (.Q(ootx_payloads_1_3), .C(clock_c), .D(n11288));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1100_1101 (.Q(ootx_payloads_1_2), .C(clock_c), .D(n11287));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1097_1098 (.Q(ootx_payloads_1_1), .C(clock_c), .D(n11286));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1094_1095 (.Q(ootx_payloads_1_0), .C(clock_c), .D(n11285));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1067_1068_adj_520 (.Q(ootx_payloads_0_263), .C(clock_c), .D(n11284));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1064_1065_adj_521 (.Q(ootx_payloads_0_262), .C(clock_c), .D(n11283));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1061_1062_adj_522 (.Q(ootx_payloads_0_261), .C(clock_c), .D(n11282));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1058_1059_adj_523 (.Q(ootx_payloads_0_260), .C(clock_c), .D(n11281));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1055_1056_adj_524 (.Q(ootx_payloads_0_259), .C(clock_c), .D(n11280));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1052_1053_adj_525 (.Q(ootx_payloads_0_258), .C(clock_c), .D(n11279));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1049_1050_adj_526 (.Q(ootx_payloads_0_257), .C(clock_c), .D(n11278));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1046_1047_adj_527 (.Q(ootx_payloads_0_256), .C(clock_c), .D(n11277));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1043_1044_adj_528 (.Q(ootx_payloads_0_255), .C(clock_c), .D(n11276));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1040_1041_adj_529 (.Q(ootx_payloads_0_254), .C(clock_c), .D(n11275));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1037_1038_adj_530 (.Q(ootx_payloads_0_253), .C(clock_c), .D(n11274));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1034_1035_adj_531 (.Q(ootx_payloads_0_252), .C(clock_c), .D(n11273));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1031_1032_adj_532 (.Q(ootx_payloads_0_251), .C(clock_c), .D(n11272));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1028_1029_adj_533 (.Q(ootx_payloads_0_250), .C(clock_c), .D(n11271));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1025_1026_adj_534 (.Q(ootx_payloads_0_249), .C(clock_c), .D(n11270));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1022_1023_adj_535 (.Q(ootx_payloads_0_248), .C(clock_c), .D(n11269));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1019_1020_adj_536 (.Q(ootx_payloads_0_247), .C(clock_c), .D(n11268));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1016_1017_adj_537 (.Q(ootx_payloads_0_246), .C(clock_c), .D(n11267));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1013_1014_adj_538 (.Q(ootx_payloads_0_245), .C(clock_c), .D(n11266));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1010_1011_adj_539 (.Q(ootx_payloads_0_244), .C(clock_c), .D(n11265));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1007_1008_adj_540 (.Q(ootx_payloads_0_243), .C(clock_c), .D(n11264));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1004_1005_adj_541 (.Q(ootx_payloads_0_242), .C(clock_c), .D(n11263));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i1001_1002_adj_542 (.Q(ootx_payloads_0_241), .C(clock_c), .D(n11262));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i998_999_adj_543 (.Q(ootx_payloads_0_240), .C(clock_c), .D(n11261));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i995_996_adj_544 (.Q(ootx_payloads_0_239), .C(clock_c), .D(n11260));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i992_993_adj_545 (.Q(ootx_payloads_0_238), .C(clock_c), .D(n11259));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i989_990_adj_546 (.Q(ootx_payloads_0_237), .C(clock_c), .D(n11258));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i986_987_adj_547 (.Q(ootx_payloads_0_236), .C(clock_c), .D(n11257));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i983_984_adj_548 (.Q(ootx_payloads_0_235), .C(clock_c), .D(n11256));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i980_981_adj_549 (.Q(ootx_payloads_0_234), .C(clock_c), .D(n11255));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i977_978_adj_550 (.Q(ootx_payloads_0_233), .C(clock_c), .D(n11254));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i974_975_adj_551 (.Q(ootx_payloads_0_232), .C(clock_c), .D(n11253));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i971_972_adj_552 (.Q(ootx_payloads_0_231), .C(clock_c), .D(n11252));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i968_969_adj_553 (.Q(ootx_payloads_0_230), .C(clock_c), .D(n11251));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i965_966_adj_554 (.Q(ootx_payloads_0_229), .C(clock_c), .D(n11250));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i962_963_adj_555 (.Q(ootx_payloads_0_228), .C(clock_c), .D(n11249));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i959_960_adj_556 (.Q(ootx_payloads_0_227), .C(clock_c), .D(n11248));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i956_957_adj_557 (.Q(ootx_payloads_0_226), .C(clock_c), .D(n11247));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i953_954_adj_558 (.Q(ootx_payloads_0_225), .C(clock_c), .D(n11246));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i950_951_adj_559 (.Q(ootx_payloads_0_224), .C(clock_c), .D(n11245));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i947_948_adj_560 (.Q(ootx_payloads_0_223), .C(clock_c), .D(n11244));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i944_945_adj_561 (.Q(ootx_payloads_0_222), .C(clock_c), .D(n11243));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i941_942_adj_562 (.Q(ootx_payloads_0_221), .C(clock_c), .D(n11242));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i938_939_adj_563 (.Q(ootx_payloads_0_220), .C(clock_c), .D(n11241));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i935_936_adj_564 (.Q(ootx_payloads_0_219), .C(clock_c), .D(n11240));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i932_933_adj_565 (.Q(ootx_payloads_0_218), .C(clock_c), .D(n11239));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i929_930_adj_566 (.Q(ootx_payloads_0_217), .C(clock_c), .D(n11238));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i926_927_adj_567 (.Q(ootx_payloads_0_216), .C(clock_c), .D(n11237));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i923_924_adj_568 (.Q(ootx_payloads_0_215), .C(clock_c), .D(n11236));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i920_921_adj_569 (.Q(ootx_payloads_0_214), .C(clock_c), .D(n11235));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i917_918_adj_570 (.Q(ootx_payloads_0_213), .C(clock_c), .D(n11234));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i914_915_adj_571 (.Q(ootx_payloads_0_212), .C(clock_c), .D(n11233));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i911_912_adj_572 (.Q(ootx_payloads_0_211), .C(clock_c), .D(n11232));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i908_909_adj_573 (.Q(ootx_payloads_0_210), .C(clock_c), .D(n11231));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i905_906_adj_574 (.Q(ootx_payloads_0_209), .C(clock_c), .D(n11230));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i902_903_adj_575 (.Q(ootx_payloads_0_208), .C(clock_c), .D(n11229));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i899_900_adj_576 (.Q(ootx_payloads_0_207), .C(clock_c), .D(n11228));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i896_897_adj_577 (.Q(ootx_payloads_0_206), .C(clock_c), .D(n11227));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i893_894_adj_578 (.Q(ootx_payloads_0_205), .C(clock_c), .D(n11226));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i890_891_adj_579 (.Q(ootx_payloads_0_204), .C(clock_c), .D(n11225));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i887_888_adj_580 (.Q(ootx_payloads_0_203), .C(clock_c), .D(n11224));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i884_885_adj_581 (.Q(ootx_payloads_0_202), .C(clock_c), .D(n11223));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i881_882_adj_582 (.Q(ootx_payloads_0_201), .C(clock_c), .D(n11222));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i878_879_adj_583 (.Q(ootx_payloads_0_200), .C(clock_c), .D(n11221));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i875_876_adj_584 (.Q(ootx_payloads_0_199), .C(clock_c), .D(n11220));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i872_873_adj_585 (.Q(ootx_payloads_0_198), .C(clock_c), .D(n11219));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i869_870_adj_586 (.Q(ootx_payloads_0_197), .C(clock_c), .D(n11218));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i866_867_adj_587 (.Q(ootx_payloads_0_196), .C(clock_c), .D(n11217));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i863_864_adj_588 (.Q(ootx_payloads_0_195), .C(clock_c), .D(n11216));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i860_861_adj_589 (.Q(ootx_payloads_0_194), .C(clock_c), .D(n11215));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i857_858_adj_590 (.Q(ootx_payloads_0_193), .C(clock_c), .D(n11214));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i854_855_adj_591 (.Q(ootx_payloads_0_192), .C(clock_c), .D(n11213));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i851_852_adj_592 (.Q(ootx_payloads_0_191), .C(clock_c), .D(n11212));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i848_849_adj_593 (.Q(ootx_payloads_0_190), .C(clock_c), .D(n11211));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i845_846_adj_594 (.Q(ootx_payloads_0_189), .C(clock_c), .D(n11210));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i842_843_adj_595 (.Q(ootx_payloads_0_188), .C(clock_c), .D(n11209));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i839_840_adj_596 (.Q(ootx_payloads_0_187), .C(clock_c), .D(n11208));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i836_837_adj_597 (.Q(ootx_payloads_0_186), .C(clock_c), .D(n11207));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i833_834_adj_598 (.Q(ootx_payloads_0_185), .C(clock_c), .D(n11206));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i830_831_adj_599 (.Q(ootx_payloads_0_184), .C(clock_c), .D(n11205));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i827_828_adj_600 (.Q(ootx_payloads_0_183), .C(clock_c), .D(n11204));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i824_825_adj_601 (.Q(ootx_payloads_0_182), .C(clock_c), .D(n11203));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i821_822_adj_602 (.Q(ootx_payloads_0_181), .C(clock_c), .D(n11202));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i818_819_adj_603 (.Q(ootx_payloads_0_180), .C(clock_c), .D(n11201));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i278_279_adj_604 (.Q(ootx_payloads_0_0), .C(clock_c), .D(n11060));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2143_12 (.CI(n22821), .I0(n3104), .I1(n3116), 
            .CO(n22822));
    SB_CARRY mod_155_add_1138_14 (.CI(n22493), .I0(n1601_adj_2150), .I1(n1631_adj_2058), 
            .CO(n22494));
    SB_LUT4 mod_155_add_1607_12_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n22617), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i815_816_adj_605 (.Q(ootx_payloads_0_179), .C(clock_c), .D(n11200));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7127_3_lut_4_lut (.I0(n954), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_216), .O(n11237));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7127_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i281_282_adj_606 (.Q(ootx_payloads_0_1), .C(clock_c), .D(n11059));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i10_3_lut (.I0(n22891), .I1(n2902), .I2(n2909), .I3(GND_net), 
            .O(n35_adj_2153));
    defparam i10_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_607 (.I0(n96), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n800));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_607.LUT_INIT = 16'h0020;
    SB_LUT4 counter_from_nskip_rise_640_add_4_23_lut (.I0(n6344), .I1(n2280), 
            .I2(counter_from_nskip_rise[21]), .I3(n22371), .O(n91[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_23_lut.LUT_INIT = 16'h8BB8;
    SB_DFF ootx_shift_registers_1_17_c (.Q(ootx_shift_registers_1_17), .C(clock_c), 
           .D(n11058));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i7641_3_lut_4_lut (.I0(n798), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1295), .O(n11751));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7641_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7049_3_lut_4_lut (.I0(n798), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_138), .O(n11159));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7049_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1138_13_lut (.I0(n1602_adj_2154), .I1(n1602_adj_2154), 
            .I2(n1631_adj_2058), .I3(n22492), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_4_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[3] ), 
            .I2(GND_net), .I3(n22307), .O(n4485[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2076_8_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n22788), .O(n3106_adj_2155)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i812_813_adj_608 (.Q(ootx_payloads_0_178), .C(clock_c), .D(n11199));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i24_4_lut (.I0(n35_adj_2153), .I1(n48_adj_2138), .I2(n44_adj_2137), 
            .I3(n36_adj_2133), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY counter_from_nskip_rise_640_add_4_23 (.CI(n22371), .I0(n2280), 
            .I1(counter_from_nskip_rise[21]), .CO(n22372));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_609 (.I0(n94_adj_1872), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n798));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_609.LUT_INIT = 16'h0020;
    SB_LUT4 i7718_3_lut_4_lut (.I0(n952), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1218), .O(n11828));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7718_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7763_3_lut_4_lut (.I0(n529), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1173), .O(n11873));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7763_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7171_3_lut_4_lut (.I0(n529), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_260), .O(n11281));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7171_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7640_3_lut_4_lut (.I0(n796), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1296), .O(n11750));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7640_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1875_7 (.CI(n22706), .I0(n2708), .I1(n2720), 
            .CO(n22707));
    SB_CARRY add_637_4 (.CI(n22307), .I0(\ootx_payloads_N_1730[3] ), .I1(GND_net), 
            .CO(n22308));
    SB_LUT4 i7048_3_lut_4_lut (.I0(n796), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_137), .O(n11158));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7048_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_18_i1_3_lut_adj_610 (.I0(bit_counters_0_18), .I1(bit_counters_1_18), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[18]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_18_i1_3_lut_adj_610.LUT_INIT = 16'hcaca;
    SB_DFF i809_810_adj_611 (.Q(ootx_payloads_0_177), .C(clock_c), .D(n11198));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i806_807_adj_612 (.Q(ootx_payloads_0_176), .C(clock_c), .D(n11197));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_10_i1_3_lut_adj_613 (.I0(bit_counters_0_26), .I1(bit_counters_1_26), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[26]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_10_i1_3_lut_adj_613.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1875_6_lut (.I0(n2709), .I1(n2709), .I2(n25192), 
            .I3(n22705), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_6_lut.LUT_INIT = 16'hA3AC;
    SB_DFF i803_804_adj_614 (.Q(ootx_payloads_0_175), .C(clock_c), .D(n11196));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i800_801_adj_615 (.Q(ootx_payloads_0_174), .C(clock_c), .D(n11195));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1607_12 (.CI(n22617), .I0(n2303), .I1(n2324), 
            .CO(n22618));
    SB_DFF i797_798_adj_616 (.Q(ootx_payloads_0_173), .C(clock_c), .D(n11194));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1607_11_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n22616), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i794_795_adj_617 (.Q(ootx_payloads_0_172), .C(clock_c), .D(n11193));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i3_4_lut_adj_618 (.I0(n2851[20]), .I1(n1212_adj_2033), .I2(n1211_adj_2031), 
            .I3(n1210_adj_2023), .O(n22873));
    defparam i3_4_lut_adj_618.LUT_INIT = 16'hfffe;
    SB_DFF i791_792_adj_619 (.Q(ootx_payloads_0_171), .C(clock_c), .D(n11192));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1138_13 (.CI(n22492), .I0(n1602_adj_2154), .I1(n1631_adj_2058), 
            .CO(n22493));
    SB_DFF i788_789_adj_620 (.Q(ootx_payloads_0_170), .C(clock_c), .D(n11191));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i785_786_adj_621 (.Q(ootx_payloads_0_169), .C(clock_c), .D(n11190));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i782_783_adj_622 (.Q(ootx_payloads_0_168), .C(clock_c), .D(n11189));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i6_4_lut_adj_623 (.I0(n1208_adj_2017), .I1(n1207_adj_2015), 
            .I2(n1204_adj_1938), .I3(n1206_adj_1980), .O(n14_adj_2156));
    defparam i6_4_lut_adj_623.LUT_INIT = 16'hfffe;
    SB_DFF i779_780_adj_624 (.Q(ootx_payloads_0_167), .C(clock_c), .D(n11188));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 counter_from_nskip_rise_640_add_4_22_lut (.I0(n6345), .I1(n2280), 
            .I2(counter_from_nskip_rise[20]), .I3(n22370), .O(n91[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_22_lut.LUT_INIT = 16'h8BB8;
    SB_DFF i776_777_adj_625 (.Q(ootx_payloads_0_166), .C(clock_c), .D(n11187));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_3_lut_adj_626 (.I0(n22873), .I1(n1202_adj_1928), .I2(n1209_adj_2021), 
            .I3(GND_net), .O(n9_adj_2157));
    defparam i1_3_lut_adj_626.LUT_INIT = 16'hecec;
    SB_LUT4 i3_4_lut_adj_627 (.I0(n2851[1]), .I1(n3112_c), .I2(n3111_adj_2158), 
            .I3(n3110_adj_2159), .O(n22889));
    defparam i3_4_lut_adj_627.LUT_INIT = 16'hfffe;
    SB_DFF i773_774_adj_628 (.Q(ootx_payloads_0_165), .C(clock_c), .D(n11186));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_629 (.I0(n82_adj_1873), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n786));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_629.LUT_INIT = 16'h0020;
    SB_DFF i770_771_adj_630 (.Q(ootx_payloads_0_164), .C(clock_c), .D(n11185));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i767_768_adj_631 (.Q(ootx_payloads_0_163), .C(clock_c), .D(n11184));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1138_12_lut (.I0(n1603), .I1(n1603), .I2(n1631_adj_2058), 
            .I3(n22491), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_637_3_lut (.I0(GND_net), .I1(\ootx_payloads_N_1730[2] ), 
            .I2(GND_net), .I3(n22306), .O(n4485[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_637_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF i764_765_adj_632 (.Q(ootx_payloads_0_162), .C(clock_c), .D(n11183));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i761_762_adj_633 (.Q(ootx_payloads_0_161), .C(clock_c), .D(n11182));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i758_759_adj_634 (.Q(ootx_payloads_0_160), .C(clock_c), .D(n11181));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_635 (.I0(n92), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n796));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_635.LUT_INIT = 16'h0020;
    SB_LUT4 i7126_3_lut_4_lut (.I0(n952), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_215), .O(n11236));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7126_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i755_756_adj_636 (.Q(ootx_payloads_0_159), .C(clock_c), .D(n11180));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i752_753_adj_637 (.Q(ootx_payloads_0_158), .C(clock_c), .D(n11179));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i749_750_adj_638 (.Q(ootx_payloads_0_157), .C(clock_c), .D(n11178));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY counter_from_nskip_rise_640_add_4_22 (.CI(n22370), .I0(n2280), 
            .I1(counter_from_nskip_rise[20]), .CO(n22371));
    SB_LUT4 i7569_3_lut_4_lut (.I0(n654), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1367), .O(n11679));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i746_747_adj_639 (.Q(ootx_payloads_0_156), .C(clock_c), .D(n11177));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7_4_lut_adj_640 (.I0(n9_adj_2157), .I1(n14_adj_2156), .I2(n1203_adj_1929), 
            .I3(n1205_adj_1940), .O(n1235_c));
    defparam i7_4_lut_adj_640.LUT_INIT = 16'hfffe;
    SB_DFF i743_744_adj_641 (.Q(ootx_payloads_0_155), .C(clock_c), .D(n11176));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1607_11 (.CI(n22616), .I0(n2304), .I1(n2324), 
            .CO(n22617));
    SB_CARRY add_637_3 (.CI(n22306), .I0(\ootx_payloads_N_1730[2] ), .I1(GND_net), 
            .CO(n22307));
    SB_DFF i740_741_adj_642 (.Q(ootx_payloads_0_154), .C(clock_c), .D(n11175));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i2_2_lut_adj_643 (.I0(n2001), .I1(n1997), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_2160));
    defparam i2_2_lut_adj_643.LUT_INIT = 16'heeee;
    SB_DFF i737_738_adj_644 (.Q(ootx_payloads_0_153), .C(clock_c), .D(n11174));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7639_3_lut_4_lut (.I0(n794), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1297), .O(n11749));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7639_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_645 (.I0(n2851[12]), .I1(n2012), .I2(n2011), 
            .I3(n2010), .O(n22942));
    defparam i3_4_lut_adj_645.LUT_INIT = 16'hfffe;
    SB_DFF i734_735_adj_646 (.Q(ootx_payloads_0_152), .C(clock_c), .D(n11173));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i11_3_lut (.I0(n22889), .I1(n3108_adj_2161), .I2(n3109_adj_2162), 
            .I3(GND_net), .O(n38_adj_2163));
    defparam i11_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7047_3_lut_4_lut (.I0(n794), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_136), .O(n11157));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7047_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7762_3_lut_4_lut (.I0(n527), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1174), .O(n11872));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7762_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i731_732_adj_647 (.Q(ootx_payloads_0_151), .C(clock_c), .D(n11172));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i728_729_adj_648 (.Q(ootx_payloads_0_150), .C(clock_c), .D(n11171));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7170_3_lut_4_lut (.I0(n527), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_259), .O(n11280));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7170_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i18_4_lut_adj_649 (.I0(n3104), .I1(n3096), .I2(n3097), .I3(n3100), 
            .O(n45_adj_2164));
    defparam i18_4_lut_adj_649.LUT_INIT = 16'hfffe;
    SB_DFF i725_726_adj_650 (.Q(ootx_payloads_0_149), .C(clock_c), .D(n11170));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1138_12 (.CI(n22491), .I0(n1603), .I1(n1631_adj_2058), 
            .CO(n22492));
    SB_LUT4 mod_155_add_1607_10_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n22615), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut_adj_651 (.I0(n2000), .I1(n2004), .I2(n1996), .I3(n2006), 
            .O(n28_adj_2165));
    defparam i12_4_lut_adj_651.LUT_INIT = 16'hfffe;
    SB_LUT4 i6977_3_lut_4_lut (.I0(n654), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_66), .O(n11087));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6977_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 counter_from_nskip_rise_640_add_4_21_lut (.I0(n6346), .I1(n2280), 
            .I2(counter_from_nskip_rise[19]), .I3(n22369), .O(n91[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_652 (.I0(n90_adj_1876), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n794));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_652.LUT_INIT = 16'h0020;
    SB_LUT4 i10_4_lut_adj_653 (.I0(n1994), .I1(n2008), .I2(n1998), .I3(n2002), 
            .O(n26_adj_2166));
    defparam i10_4_lut_adj_653.LUT_INIT = 16'hfffe;
    SB_LUT4 i7638_3_lut_4_lut (.I0(n792), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1298), .O(n11748));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7638_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7046_3_lut_4_lut (.I0(n792), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_135), .O(n11156));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7046_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i722_723_adj_654 (.Q(ootx_payloads_0_148), .C(clock_c), .D(n11169));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i11_4_lut_adj_655 (.I0(n1999), .I1(n2007), .I2(n2005), .I3(n2003), 
            .O(n27_adj_2167));
    defparam i11_4_lut_adj_655.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_656 (.I0(n3102), .I1(n3086), .I2(n3107_adj_2168), 
            .I3(n3089), .O(n42_adj_2169));
    defparam i15_4_lut_adj_656.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_657 (.I0(n22942), .I1(n18_adj_2160), .I2(n1995), 
            .I3(n2009), .O(n25_adj_2170));
    defparam i9_4_lut_adj_657.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_658 (.I0(n25_adj_2170), .I1(n27_adj_2167), .I2(n26_adj_2166), 
            .I3(n28_adj_2165), .O(n2027));
    defparam i15_4_lut_adj_658.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1875_6 (.CI(n22705), .I0(n2709), .I1(n25192), 
            .CO(n22706));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_659 (.I0(n80), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n784));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_659.LUT_INIT = 16'h0020;
    SB_LUT4 i7717_3_lut_4_lut (.I0(n950), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1219), .O(n11827));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7717_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2143_11_lut (.I0(n3105_adj_2136), .I1(n3105_adj_2136), 
            .I2(n3116), .I3(n22820), .O(n19_adj_1967)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1138_11_lut (.I0(n1604), .I1(n1604), .I2(n1631_adj_2058), 
            .I3(n22490), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7637_3_lut_4_lut (.I0(n790), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1299), .O(n11747));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7637_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_637_2 (.CI(GND_net), .I0(\ootx_payloads_N_1730[1] ), .I1(\ootx_payloads_N_1730[1] ), 
            .CO(n22306));
    SB_CARRY counter_from_nskip_rise_640_add_4_21 (.CI(n22369), .I0(n2280), 
            .I1(counter_from_nskip_rise[19]), .CO(n22370));
    SB_LUT4 i7045_3_lut_4_lut (.I0(n790), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_134), .O(n11155));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7045_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_9_i1_3_lut_adj_660 (.I0(bit_counters_0_27), .I1(bit_counters_1_27), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[27]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_9_i1_3_lut_adj_660.LUT_INIT = 16'hcaca;
    SB_LUT4 i7761_3_lut_4_lut (.I0(n525), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1175), .O(n11871));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7761_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_2_lut (.I0(n3090), .I1(n3083), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_2171));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7169_3_lut_4_lut (.I0(n525), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_258), .O(n11279));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7169_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19415_2_lut_4_lut (.I0(n19_adj_2172), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24065));
    defparam i19415_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_LUT4 i7125_3_lut_4_lut (.I0(n950), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_214), .O(n11235));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7125_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19430_2_lut_4_lut (.I0(n19_adj_2172), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24095));
    defparam i19430_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 i7636_3_lut_4_lut (.I0(n788), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1300), .O(n11746));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7636_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7044_3_lut_4_lut (.I0(n788), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_133), .O(n11154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7044_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7635_3_lut_4_lut (.I0(n786), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1301), .O(n11745));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7635_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1942_28 (.CI(n22753), .I0(n2787), .I1(n2819), 
            .CO(n22754));
    SB_LUT4 i7043_3_lut_4_lut (.I0(n786), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_132), .O(n11153));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7043_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_355_33_lut (.I0(GND_net), .I1(\counter_from_last_rise[31] ), 
            .I2(GND_net), .I3(n22305), .O(n6334)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_661 (.I0(n78_adj_1891), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n782));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_661.LUT_INIT = 16'h0020;
    SB_LUT4 mod_155_add_1875_5_lut (.I0(n2710), .I1(n2710), .I2(n2720), 
            .I3(n22704), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_27_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n22752), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7634_3_lut_4_lut (.I0(n784), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1302), .O(n11744));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7634_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7042_3_lut_4_lut (.I0(n784), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_131), .O(n11152));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7042_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7568_3_lut_4_lut (.I0(n652), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1368), .O(n11678));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i18_2_lut_3_lut (.I0(n6_adj_2054), .I1(ootx_payloads_N_1699[1]), 
            .I2(ootx_payloads_N_1699[2]), .I3(GND_net), .O(n18_adj_2173));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(119[37:62])
    defparam EnabledDecoder_2_i18_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i19_2_lut_3_lut (.I0(n6_adj_2054), .I1(ootx_payloads_N_1699[1]), 
            .I2(ootx_payloads_N_1699[2]), .I3(GND_net), .O(n19_adj_2172));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(119[37:62])
    defparam EnabledDecoder_2_i19_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i7760_3_lut_4_lut (.I0(n523), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1176), .O(n11870));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7760_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6976_3_lut_4_lut (.I0(n652), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_65), .O(n11086));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7168_3_lut_4_lut (.I0(n523), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_257), .O(n11278));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7168_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7633_3_lut_4_lut (.I0(n782), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1303), .O(n11743));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7633_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut_adj_662 (.I0(n3106_adj_2155), .I1(n3091), .I2(n3095), 
            .I3(n3103), .O(n44_adj_2174));
    defparam i17_4_lut_adj_662.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1607_10 (.CI(n22615), .I0(n2305), .I1(n2324), 
            .CO(n22616));
    SB_LUT4 i7041_3_lut_4_lut (.I0(n782), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_130), .O(n11151));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7041_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_1875_5 (.CI(n22704), .I0(n2710), .I1(n2720), 
            .CO(n22705));
    SB_CARRY mod_155_add_2143_11 (.CI(n22820), .I0(n3105_adj_2136), .I1(n3116), 
            .CO(n22821));
    SB_LUT4 i23_4_lut_adj_663 (.I0(n45_adj_2164), .I1(n3087), .I2(n38_adj_2163), 
            .I3(n3092), .O(n50_adj_2175));
    defparam i23_4_lut_adj_663.LUT_INIT = 16'hfffe;
    SB_LUT4 i7716_3_lut_4_lut (.I0(n948), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1220), .O(n11826));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7716_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7632_3_lut_4_lut (.I0(n780), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1304), .O(n11742));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7040_3_lut_4_lut (.I0(n780), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_129), .O(n11150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7040_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i21_4_lut_adj_664 (.I0(n3094), .I1(n42_adj_2169), .I2(n3093), 
            .I3(n3099), .O(n48_adj_2177));
    defparam i21_4_lut_adj_664.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1138_11 (.CI(n22490), .I0(n1604), .I1(n1631_adj_2058), 
            .CO(n22491));
    SB_LUT4 mod_155_add_1607_9_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n22614), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_665 (.I0(n76), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n780));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_665.LUT_INIT = 16'h0020;
    SB_LUT4 i7631_3_lut_4_lut (.I0(n778), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1305), .O(n11741));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7631_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22_4_lut_adj_666 (.I0(n3084), .I1(n44_adj_2174), .I2(n32_adj_2171), 
            .I3(n3088), .O(n49_adj_2179));
    defparam i22_4_lut_adj_666.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1607_9 (.CI(n22614), .I0(n2306), .I1(n2324), 
            .CO(n22615));
    SB_LUT4 i7039_3_lut_4_lut (.I0(n778), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_128), .O(n11149));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7039_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7124_3_lut_4_lut (.I0(n948), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_213), .O(n11234));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7124_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19414_2_lut_4_lut (.I0(n12_adj_2180), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24063));
    defparam i19414_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_LUT4 i19429_2_lut_4_lut (.I0(n12_adj_2180), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24093));
    defparam i19429_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 i20_4_lut_adj_667 (.I0(n3098), .I1(n3085), .I2(n3101), .I3(n3105_adj_2136), 
            .O(n47_adj_2181));
    defparam i20_4_lut_adj_667.LUT_INIT = 16'hfffe;
    SB_LUT4 counter_from_nskip_rise_640_add_4_20_lut (.I0(n6333[18]), .I1(n2280), 
            .I2(counter_from_nskip_rise[18]), .I3(n22368), .O(n91[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i7715_3_lut_4_lut (.I0(n946), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1221), .O(n11825));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7715_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i26_4_lut_adj_668 (.I0(n47_adj_2181), .I1(n49_adj_2179), .I2(n48_adj_2177), 
            .I3(n50_adj_2175), .O(n3116));
    defparam i26_4_lut_adj_668.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1138_10_lut (.I0(n1605), .I1(n1605), .I2(n1631_adj_2058), 
            .I3(n22489), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20513_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25181));
    defparam i20513_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_355_32_lut (.I0(GND_net), .I1(\counter_from_last_rise[30] ), 
            .I2(GND_net), .I3(n22304), .O(n6335)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut_4_lut_adj_669 (.I0(n11_adj_2039), 
            .I1(ootx_payloads_N_1699[1]), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(ootx_payloads_N_1699[2]), .O(n39_adj_1902));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i39_2_lut_3_lut_4_lut_adj_669.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut_adj_670 (.I0(n11_adj_2039), 
            .I1(ootx_payloads_N_1699[1]), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(ootx_payloads_N_1699[2]), .O(n40_adj_2049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut_adj_670.LUT_INIT = 16'h0800;
    SB_LUT4 i4_2_lut_adj_671 (.I0(n2589), .I1(n2608), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_2182));
    defparam i4_2_lut_adj_671.LUT_INIT = 16'heeee;
    SB_LUT4 i7759_3_lut_4_lut (.I0(n521), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1177), .O(n11869));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7759_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7123_3_lut_4_lut (.I0(n946), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_212), .O(n11233));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7123_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY mod_155_add_2076_8 (.CI(n22788), .I0(n3007), .I1(n3017), 
            .CO(n22789));
    SB_LUT4 i7167_3_lut_4_lut (.I0(n521), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_256), .O(n11277));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7167_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_20 (.CI(n22368), .I0(n2280), 
            .I1(counter_from_nskip_rise[18]), .CO(n22369));
    SB_LUT4 i14_4_lut_adj_672 (.I0(n2601), .I1(n2592), .I2(n2605), .I3(n2588), 
            .O(n36_adj_2183));
    defparam i14_4_lut_adj_672.LUT_INIT = 16'hfffe;
    SB_LUT4 i7567_3_lut_4_lut (.I0(n650), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1369), .O(n11677));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2143_10_lut (.I0(n3106_adj_2155), .I1(n3106_adj_2155), 
            .I2(n3116), .I3(n22819), .O(n17_adj_1965)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7630_3_lut_4_lut (.I0(n776), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1306), .O(n11740));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7630_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7038_3_lut_4_lut (.I0(n776), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_127), .O(n11148));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7038_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_673 (.I0(n2851[6]), .I1(n2612), .I2(n2611), .I3(n2610), 
            .O(n22894));
    defparam i3_4_lut_adj_673.LUT_INIT = 16'hfffe;
    SB_LUT4 i7629_3_lut_4_lut (.I0(n774), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1307), .O(n11739));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7629_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_adj_674 (.I0(n2603), .I1(n2606), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_2184));
    defparam i2_2_lut_adj_674.LUT_INIT = 16'heeee;
    SB_LUT4 i7037_3_lut_4_lut (.I0(n774), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_126), .O(n11147));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7037_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_1607_8_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n22613), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_32 (.CI(n22304), .I0(\counter_from_last_rise[30] ), 
            .I1(GND_net), .CO(n22305));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_675 (.I0(n74_adj_1899), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n778));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_675.LUT_INIT = 16'h0020;
    SB_LUT4 i6975_3_lut_4_lut (.I0(n650), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_64), .O(n11085));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6975_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF ootx_shift_registers_1_16_c (.Q(ootx_shift_registers_1_16), .C(clock_c), 
           .D(n11057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i19413_2_lut_4_lut (.I0(n14_adj_2149), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24061));
    defparam i19413_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_LUT4 i7714_3_lut_4_lut (.I0(n944), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1222), .O(n11824));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7714_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19428_2_lut_4_lut (.I0(n14_adj_2149), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24091));
    defparam i19428_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 i7009_3_lut_4_lut (.I0(n718), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_98), .O(n11119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7009_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7601_3_lut_4_lut (.I0(n718), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1335), .O(n11711));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7601_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_adj_676 (.I0(n22894), .I1(n2596), .I2(n2609), .I3(GND_net), 
            .O(n23_adj_2185));
    defparam i1_3_lut_adj_676.LUT_INIT = 16'hecec;
    SB_LUT4 i7758_3_lut_4_lut (.I0(n1032), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1178), .O(n11868));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7758_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7166_3_lut_4_lut (.I0(n1032), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_255), .O(n11276));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7166_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_677 (.I0(n77), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n974));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_677.LUT_INIT = 16'h0080;
    SB_LUT4 i18_4_lut_adj_678 (.I0(n2599), .I1(n36_adj_2183), .I2(n26_adj_2182), 
            .I3(n2598), .O(n40_adj_2186));
    defparam i18_4_lut_adj_678.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1138_10 (.CI(n22489), .I0(n1605), .I1(n1631_adj_2058), 
            .CO(n22490));
    SB_CARRY mod_155_add_1607_8 (.CI(n22613), .I0(n2307), .I1(n2324), 
            .CO(n22614));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_679 (.I0(n135), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n1032));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_679.LUT_INIT = 16'h0080;
    SB_LUT4 counter_from_nskip_rise_640_add_4_19_lut (.I0(n6333[17]), .I1(n2280), 
            .I2(counter_from_nskip_rise[17]), .I3(n22367), .O(n91[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i7122_3_lut_4_lut (.I0(n944), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_211), .O(n11232));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7122_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_8_i1_3_lut_adj_680 (.I0(bit_counters_0_28), .I1(bit_counters_1_28), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[28]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_8_i1_3_lut_adj_680.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1138_9_lut (.I0(n1606), .I1(n1606), .I2(n1631_adj_2058), 
            .I3(n22488), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_681 (.I0(n2595), .I1(n2590), .I2(n2604), .I3(n2602), 
            .O(n38_adj_2187));
    defparam i16_4_lut_adj_681.LUT_INIT = 16'hfffe;
    SB_LUT4 EnabledDecoder_2_i78_2_lut_3_lut (.I0(n30_adj_1855), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n78_adj_1891));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i78_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i17_4_lut_adj_682 (.I0(n2600), .I1(n23_adj_2185), .I2(n2597), 
            .I3(n24_adj_2184), .O(n39_adj_2188));
    defparam i17_4_lut_adj_682.LUT_INIT = 16'hfffe;
    SB_LUT4 EnabledDecoder_2_i77_2_lut_3_lut (.I0(n30_adj_1855), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n77));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i77_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i15_4_lut_adj_683 (.I0(n2593), .I1(n2594), .I2(n2591), .I3(n2607), 
            .O(n37_adj_2189));
    defparam i15_4_lut_adj_683.LUT_INIT = 16'hfffe;
    SB_CARRY counter_from_nskip_rise_640_add_4_19 (.CI(n22367), .I0(n2280), 
            .I1(counter_from_nskip_rise[17]), .CO(n22368));
    SB_LUT4 Mux_7_i1_3_lut (.I0(bit_counters_0_29), .I1(bit_counters_1_29), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[29]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_7_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_355_31_lut (.I0(GND_net), .I1(\counter_from_last_rise[29] ), 
            .I2(GND_net), .I3(n22303), .O(n6336)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_4_lut_adj_684 (.I0(n37_adj_2189), .I1(n39_adj_2188), .I2(n38_adj_2187), 
            .I3(n40_adj_2186), .O(n2621));
    defparam i21_4_lut_adj_684.LUT_INIT = 16'hfffe;
    SB_LUT4 Mux_6_i1_3_lut (.I0(bit_counters_0_30), .I1(bit_counters_1_30), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[30]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_6_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_2_lut (.I0(n2792), .I1(n2790), .I2(GND_net), .I3(GND_net), 
            .O(n30_adj_2190));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_155_add_1875_4_lut (.I0(n2711), .I1(n2711), .I2(n2720), 
            .I3(n22703), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_31 (.CI(n22303), .I0(\counter_from_last_rise[29] ), 
            .I1(GND_net), .CO(n22304));
    SB_LUT4 i16_4_lut_adj_685 (.I0(n2795), .I1(n2807), .I2(n2797), .I3(n2806), 
            .O(n40_adj_2191));
    defparam i16_4_lut_adj_685.LUT_INIT = 16'hfffe;
    SB_LUT4 i7564_3_lut_4_lut (.I0(n644), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1372), .O(n11674));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2076_7_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n22787), .O(n3107_adj_2168)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1607_7_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n22612), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF ootx_shift_registers_1_15_c (.Q(ootx_shift_registers_1_15), .C(clock_c), 
           .D(n11056));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_CARRY mod_155_add_1875_4 (.CI(n22703), .I0(n2711), .I1(n2720), 
            .CO(n22704));
    SB_LUT4 i3_4_lut_adj_686 (.I0(n2851[4]), .I1(n2812), .I2(n2811), .I3(n2810), 
            .O(n22892));
    defparam i3_4_lut_adj_686.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_687 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n162_adj_1905), .I3(GND_net), .O(n802));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_687.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_688 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n164), .I3(GND_net), .O(n804));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_688.LUT_INIT = 16'h4040;
    SB_LUT4 i14_4_lut_adj_689 (.I0(n2789), .I1(n2798), .I2(n2808), .I3(n2804), 
            .O(n38_adj_2192));
    defparam i14_4_lut_adj_689.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_690 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n166_adj_2018), .I3(GND_net), .O(n806));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_690.LUT_INIT = 16'h4040;
    SB_LUT4 i1_3_lut_adj_691 (.I0(n2788), .I1(n22892), .I2(n2809), .I3(GND_net), 
            .O(n25_adj_2193));
    defparam i1_3_lut_adj_691.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_3_lut_adj_692 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n168), .I3(GND_net), .O(n808));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_692.LUT_INIT = 16'h4040;
    SB_LUT4 i20_4_lut_adj_693 (.I0(n2799), .I1(n40_adj_2191), .I2(n30_adj_2190), 
            .I3(n2796), .O(n44_adj_2194));
    defparam i20_4_lut_adj_693.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1138_9 (.CI(n22488), .I0(n1606), .I1(n1631_adj_2058), 
            .CO(n22489));
    SB_CARRY mod_155_add_1607_7 (.CI(n22612), .I0(n2308), .I1(n2324), 
            .CO(n22613));
    SB_LUT4 i1_2_lut_3_lut_adj_694 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n170_adj_2042), .I3(GND_net), .O(n810));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_694.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_695 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n172), .I3(GND_net), .O(n812));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_695.LUT_INIT = 16'h4040;
    SB_LUT4 counter_from_nskip_rise_640_add_4_18_lut (.I0(n6333[16]), .I1(n2280), 
            .I2(counter_from_nskip_rise[16]), .I3(n22366), .O(n91[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_18_lut.LUT_INIT = 16'h8BB8;
    SB_DFF ootx_shift_registers_1_14_c (.Q(ootx_shift_registers_1_14), .C(clock_c), 
           .D(n11055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i18_4_lut_adj_696 (.I0(n2802), .I1(n2793), .I2(n2805), .I3(n2803), 
            .O(n42_adj_2195));
    defparam i18_4_lut_adj_696.LUT_INIT = 16'hfffe;
    SB_LUT4 EnabledDecoder_2_i113_2_lut_4_lut (.I0(n17_adj_1864), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n113));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i113_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY mod_155_add_2143_10 (.CI(n22819), .I0(n3106_adj_2155), .I1(n3116), 
            .CO(n22820));
    SB_LUT4 mod_155_add_1138_8_lut (.I0(n1607), .I1(n1607), .I2(n1631_adj_2058), 
            .I3(n22487), .O(n1706_adj_1810)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_355_30_lut (.I0(GND_net), .I1(\counter_from_last_rise[28] ), 
            .I2(GND_net), .I3(n22302), .O(n6337)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_from_nskip_rise_640_add_4_18 (.CI(n22366), .I0(n2280), 
            .I1(counter_from_nskip_rise[16]), .CO(n22367));
    SB_LUT4 mod_155_add_1607_6_lut (.I0(n2309), .I1(n2309), .I2(n25198), 
            .I3(n22611), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_6_lut.LUT_INIT = 16'hA3AC;
    SB_DFF ootx_shift_registers_1_13_c (.Q(ootx_shift_registers_1_13), .C(clock_c), 
           .D(n11054));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_CARRY mod_155_add_1138_8 (.CI(n22487), .I0(n1607), .I1(n1631_adj_2058), 
            .CO(n22488));
    SB_CARRY add_355_30 (.CI(n22302), .I0(\counter_from_last_rise[28] ), 
            .I1(GND_net), .CO(n22303));
    SB_LUT4 EnabledDecoder_2_i111_2_lut_4_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n111));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i111_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i19_4_lut_adj_697 (.I0(n25_adj_2193), .I1(n38_adj_2192), .I2(n2794), 
            .I3(n2801), .O(n43_adj_2196));
    defparam i19_4_lut_adj_697.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1607_6 (.CI(n22611), .I0(n2309), .I1(n25198), 
            .CO(n22612));
    SB_DFF ootx_shift_registers_1_12_c (.Q(ootx_shift_registers_1_12), .C(clock_c), 
           .D(n11053));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_698 (.I0(ootx_payloads_N_1744[1]), .I1(ootx_payloads_N_1744[0]), 
            .I2(new_data), .I3(reset_c), .O(n9513));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_3_lut_4_lut_adj_698.LUT_INIT = 16'h00e0;
    SB_LUT4 counter_from_nskip_rise_640_add_4_17_lut (.I0(n6333[15]), .I1(n2280), 
            .I2(counter_from_nskip_rise[15]), .I3(n22365), .O(n91[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_adj_699 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n218), .I3(GND_net), .O(n858));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_699.LUT_INIT = 16'h4040;
    SB_LUT4 Mux_23_i1_3_lut_adj_700 (.I0(bit_counters_0_13), .I1(bit_counters_1_13), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[13]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_23_i1_3_lut_adj_700.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_4_lut_adj_701 (.I0(n2800), .I1(n2786), .I2(n2791), .I3(n2787), 
            .O(n41_adj_2197));
    defparam i17_4_lut_adj_701.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1138_7_lut (.I0(n1608), .I1(n1608), .I2(n1631_adj_2058), 
            .I3(n22486), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_adj_702 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n220), .I3(GND_net), .O(n860));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_702.LUT_INIT = 16'h4040;
    SB_LUT4 add_355_29_lut (.I0(GND_net), .I1(\counter_from_last_rise[27] ), 
            .I2(GND_net), .I3(n22301), .O(n6338)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23_4_lut_adj_703 (.I0(n41_adj_2197), .I1(n43_adj_2196), .I2(n42_adj_2195), 
            .I3(n44_adj_2194), .O(n2819));
    defparam i23_4_lut_adj_703.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_704 (.I0(ootx_payloads_N_1698), .I1(ootx_payloads_N_1744[0]), 
            .I2(ootx_payloads_N_1744[1]), .I3(\lighthouse[0] ), .O(n22943));
    defparam i2_3_lut_4_lut_adj_704.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_705 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n226), .I3(GND_net), .O(n866));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_705.LUT_INIT = 16'h4040;
    SB_CARRY counter_from_nskip_rise_640_add_4_17 (.CI(n22365), .I0(n2280), 
            .I1(counter_from_nskip_rise[15]), .CO(n22366));
    SB_LUT4 i2_2_lut_adj_706 (.I0(n1512), .I1(n1510), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_2198));
    defparam i2_2_lut_adj_706.LUT_INIT = 16'heeee;
    SB_CARRY mod_155_add_2076_7 (.CI(n22787), .I0(n3008), .I1(n3017), 
            .CO(n22788));
    SB_LUT4 i1_2_lut_3_lut_adj_707 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n234), .I3(GND_net), .O(n874));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_707.LUT_INIT = 16'h4040;
    SB_CARRY add_355_29 (.CI(n22301), .I0(\counter_from_last_rise[27] ), 
            .I1(GND_net), .CO(n22302));
    SB_DFF ootx_shift_registers_1_11_c (.Q(ootx_shift_registers_1_11), .C(clock_c), 
           .D(n11052));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i15352_4_lut (.I0(n2851[17]), .I1(n1509), .I2(n6_adj_2198), 
            .I3(n1511), .O(n19448));
    defparam i15352_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i7_4_lut_adj_708 (.I0(n1505), .I1(n1504), .I2(n1506), .I3(n19448), 
            .O(n18_adj_2199));
    defparam i7_4_lut_adj_708.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1942_27 (.CI(n22752), .I0(n2788), .I1(n2819), 
            .CO(n22753));
    SB_LUT4 mod_155_add_2076_6_lut (.I0(n3009), .I1(n3009), .I2(n25183), 
            .I3(n22786), .O(n3108_adj_2161)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_155_add_2143_9_lut (.I0(n3107_adj_2168), .I1(n3107_adj_2168), 
            .I2(n3116), .I3(n22818), .O(n15_adj_1955)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1875_3_lut (.I0(n2712), .I1(n2712), .I2(n2720), 
            .I3(n22702), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_3_lut.LUT_INIT = 16'hCA3A;
    SB_DFF ootx_shift_registers_1_10_c (.Q(ootx_shift_registers_1_10), .C(clock_c), 
           .D(n11051));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_adj_709 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n250), .I3(GND_net), .O(n890));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_709.LUT_INIT = 16'h4040;
    SB_CARRY mod_155_add_2076_6 (.CI(n22786), .I0(n3009), .I1(n25183), 
            .CO(n22787));
    SB_LUT4 i5_2_lut_adj_710 (.I0(n1503), .I1(n1502), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_2200));
    defparam i5_2_lut_adj_710.LUT_INIT = 16'heeee;
    SB_DFF ootx_shift_registers_1_9_c (.Q(ootx_shift_registers_1_9), .C(clock_c), 
           .D(n11050));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i9_4_lut_adj_711 (.I0(n1508), .I1(n18_adj_2199), .I2(n1507), 
            .I3(n1501), .O(n20_adj_2201));
    defparam i9_4_lut_adj_711.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_712 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n252), .I3(GND_net), .O(n892));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_712.LUT_INIT = 16'h4040;
    SB_DFF ootx_shift_registers_1_8_c (.Q(ootx_shift_registers_1_8), .C(clock_c), 
           .D(n11049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_adj_713 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n256), .I3(GND_net), .O(n896));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_713.LUT_INIT = 16'h4040;
    SB_LUT4 mod_155_add_1607_5_lut (.I0(n2310), .I1(n2310), .I2(n2324), 
            .I3(n22610), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1942_26_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n22751), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut_adj_714 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n258), .I3(GND_net), .O(n898));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_714.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_715 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n260), .I3(GND_net), .O(n900));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_715.LUT_INIT = 16'h4040;
    SB_LUT4 i10_4_lut_adj_716 (.I0(n1499), .I1(n20_adj_2201), .I2(n16_adj_2200), 
            .I3(n1500), .O(n1532));
    defparam i10_4_lut_adj_716.LUT_INIT = 16'hfffe;
    SB_DFF ootx_shift_registers_1_7_c (.Q(ootx_shift_registers_1_7), .C(clock_c), 
           .D(n11048));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_adj_717 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n262), .I3(GND_net), .O(n902));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_717.LUT_INIT = 16'h4040;
    SB_DFF ootx_shift_registers_1_6_c (.Q(ootx_shift_registers_1_6), .C(clock_c), 
           .D(n11047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i6692_2_lut (.I0(data), .I1(ootx_payloads_N_1744[0]), .I2(GND_net), 
            .I3(GND_net), .O(n10802));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[6] 189[13])
    defparam i6692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_718 (.I0(new_data), .I1(\lighthouse[0] ), .I2(n25222), 
            .I3(GND_net), .O(n23147));
    defparam i1_3_lut_adj_718.LUT_INIT = 16'h8080;
    SB_DFF ootx_shift_registers_1_5_c (.Q(ootx_shift_registers_1_5), .C(clock_c), 
           .D(n11046));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 mux_430_Mux_1_i3_4_lut (.I0(n10802), .I1(n30), .I2(ootx_payloads_N_1744[1]), 
            .I3(\lighthouse[0] ), .O(ootx_states_1__1__N_896[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[6] 189[13])
    defparam mux_430_Mux_1_i3_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 Mux_23_i1_3_lut_adj_719 (.I0(data_counters_0_15), .I1(data_counters_1_15), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1699[15] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(172[25:35])
    defparam Mux_23_i1_3_lut_adj_719.LUT_INIT = 16'hcaca;
    SB_DFF ootx_shift_registers_1_4_c (.Q(ootx_shift_registers_1_4), .C(clock_c), 
           .D(n11045));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFF i719_720_adj_720 (.Q(ootx_payloads_0_147), .C(clock_c), .D(n11168));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_8_i1_3_lut_adj_721 (.I0(payload_lengths_0_12), .I1(payload_lengths_1_12), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[12] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_8_i1_3_lut_adj_721.LUT_INIT = 16'hcaca;
    SB_DFF ootx_shift_registers_1_3_c (.Q(ootx_shift_registers_1_3), .C(clock_c), 
           .D(n11044));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFF ootx_shift_registers_1_2_c (.Q(ootx_shift_registers_1_2), .C(clock_c), 
           .D(n11043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFF ootx_shift_registers_1_1_c (.Q(ootx_shift_registers_1_1), .C(clock_c), 
           .D(n11042));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 Mux_36_i1_3_lut_adj_722 (.I0(bit_counters_0_0), .I1(bit_counters_1_0), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_36_i1_3_lut_adj_722.LUT_INIT = 16'hcaca;
    SB_DFF ootx_shift_registers_1_0_c (.Q(ootx_shift_registers_1_0), .C(clock_c), 
           .D(n11041));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_CARRY mod_155_add_1138_7 (.CI(n22486), .I0(n1608), .I1(n1631_adj_2058), 
            .CO(n22487));
    SB_DFF ootx_shift_registers_0_17_c (.Q(ootx_shift_registers_0_17), .C(clock_c), 
           .D(n11040));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 Mux_20_i1_3_lut_adj_723 (.I0(payload_lengths_0_0), .I1(payload_lengths_1_0), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[0] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_20_i1_3_lut_adj_723.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_35_i1_3_lut_adj_724 (.I0(bit_counters_0_1), .I1(bit_counters_1_1), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_35_i1_3_lut_adj_724.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_from_nskip_rise_640_add_4_16_lut (.I0(n6333[14]), .I1(n2280), 
            .I2(counter_from_nskip_rise[14]), .I3(n22364), .O(n91[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_16_lut.LUT_INIT = 16'h8BB8;
    SB_DFF ootx_shift_registers_0_16_c (.Q(ootx_shift_registers_0_16), .C(clock_c), 
           .D(n11039));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 Mux_34_i1_3_lut_adj_725 (.I0(bit_counters_0_2), .I1(bit_counters_1_2), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[2]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_34_i1_3_lut_adj_725.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1138_6_lut (.I0(n1609), .I1(n1609), .I2(n25199), 
            .I3(n22485), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i20518_1_lut (.I0(n1334_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25186));
    defparam i20518_1_lut.LUT_INIT = 16'h5555;
    SB_DFF ootx_shift_registers_0_15_c (.Q(ootx_shift_registers_0_15), .C(clock_c), 
           .D(n11038));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_adj_726 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n161), .I3(GND_net), .O(n930));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_726.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_727 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n163), .I3(GND_net), .O(n932));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_727.LUT_INIT = 16'h4040;
    SB_CARRY counter_from_nskip_rise_640_add_4_16 (.CI(n22364), .I0(n2280), 
            .I1(counter_from_nskip_rise[14]), .CO(n22365));
    SB_CARRY mod_155_add_1875_3 (.CI(n22702), .I0(n2712), .I1(n2720), 
            .CO(n22703));
    SB_CARRY mod_155_add_1607_5 (.CI(n22610), .I0(n2310), .I1(n2324), 
            .CO(n22611));
    SB_LUT4 i1_2_lut_3_lut_adj_728 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n165), .I3(GND_net), .O(n934));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_728.LUT_INIT = 16'h4040;
    SB_DFFESR sensor_state_switch_counter_641__i5 (.Q(sensor_state_switch_counter[5]), 
            .C(clock_c), .E(n13338), .D(n100[5]), .R(n13346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    SB_LUT4 i20517_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25185));
    defparam i20517_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_729 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n167), .I3(GND_net), .O(n936));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_729.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_730 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n169), .I3(GND_net), .O(n938));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_730.LUT_INIT = 16'h4040;
    SB_DFF ootx_shift_registers_0_14_c (.Q(ootx_shift_registers_0_14), .C(clock_c), 
           .D(n11037));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_adj_731 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n171), .I3(GND_net), .O(n940));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_731.LUT_INIT = 16'h4040;
    SB_DFFESR sensor_state_switch_counter_641__i4 (.Q(sensor_state_switch_counter[4]), 
            .C(clock_c), .E(n13338), .D(n100[4]), .R(n13346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    SB_DFFESR sensor_state_switch_counter_641__i3 (.Q(sensor_state_switch_counter[3]), 
            .C(clock_c), .E(n13338), .D(n100[3]), .R(n13346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    SB_DFF ootx_shift_registers_0_13_c (.Q(ootx_shift_registers_0_13), .C(clock_c), 
           .D(n11036));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFFESR sensor_state_switch_counter_641__i2 (.Q(sensor_state_switch_counter[2]), 
            .C(clock_c), .E(n13338), .D(n100[2]), .R(n13346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    SB_DFFESR sensor_state_switch_counter_641__i1 (.Q(sensor_state_switch_counter[1]), 
            .C(clock_c), .E(n13338), .D(n100[1]), .R(n13346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    SB_DFF ootx_shift_registers_0_12_c (.Q(ootx_shift_registers_0_12), .C(clock_c), 
           .D(n11035));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFFESR sync__i1 (.Q(sync[1]), .C(clock_c), .E(n2282), .D(n20098), 
            .R(n18844));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_DFF ootx_shift_registers_0_11_c (.Q(ootx_shift_registers_0_11), .C(clock_c), 
           .D(n11034));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 EnabledDecoder_2_i116_2_lut_3_lut (.I0(n36_adj_2041), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n116));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i116_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF ootx_shift_registers_0_10_c (.Q(ootx_shift_registers_0_10), .C(clock_c), 
           .D(n11033));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 Mux_19_i1_3_lut_adj_732 (.I0(bit_counters_0_17), .I1(bit_counters_1_17), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[17]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_19_i1_3_lut_adj_732.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_155_add_1607_4_lut (.I0(n2311), .I1(n2311), .I2(n2324), 
            .I3(n22609), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF ootx_shift_registers_0_9_c (.Q(ootx_shift_registers_0_9), .C(clock_c), 
           .D(n11032));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 add_355_28_lut (.I0(GND_net), .I1(\counter_from_last_rise[26] ), 
            .I2(GND_net), .I3(n22300), .O(n6339)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_2076_5_lut (.I0(n3010), .I1(n3010), .I2(n3017), 
            .I3(n22785), .O(n3109_adj_2162)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF ootx_shift_registers_0_8_c (.Q(ootx_shift_registers_0_8), .C(clock_c), 
           .D(n11031));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFF ootx_shift_registers_0_7_c (.Q(ootx_shift_registers_0_7), .C(clock_c), 
           .D(n11030));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_CARRY mod_155_add_1138_6 (.CI(n22485), .I0(n1609), .I1(n25199), 
            .CO(n22486));
    SB_DFF ootx_shift_registers_0_6_c (.Q(ootx_shift_registers_0_6), .C(clock_c), 
           .D(n11029));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_733 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n125), .O(n1022));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_733.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_734 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n93_adj_2014), .O(n990));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_734.LUT_INIT = 16'h4000;
    SB_DFF ootx_shift_registers_0_5_c (.Q(ootx_shift_registers_0_5), .C(clock_c), 
           .D(n11028));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 EnabledDecoder_2_i115_2_lut_3_lut (.I0(n36_adj_2041), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n115));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i115_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_735 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n115), .O(n1012));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_735.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_736 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n117), .O(n1014));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_736.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_737 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n136), .O(n968));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_737.LUT_INIT = 16'h4000;
    SB_LUT4 counter_from_nskip_rise_640_add_4_15_lut (.I0(n6333[13]), .I1(n2280), 
            .I2(counter_from_nskip_rise[13]), .I3(n22363), .O(n91[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_15_lut.LUT_INIT = 16'h8BB8;
    SB_DFF ootx_shift_registers_0_4_c (.Q(ootx_shift_registers_0_4), .C(clock_c), 
           .D(n11027));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_738 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n87), .O(n984));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_738.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_739 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n73), .O(n970));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_739.LUT_INIT = 16'h4000;
    SB_CARRY add_355_28 (.CI(n22300), .I0(\counter_from_last_rise[26] ), 
            .I1(GND_net), .CO(n22301));
    SB_LUT4 EnabledDecoder_2_i107_2_lut (.I0(n43_adj_1944), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i107_2_lut.LUT_INIT = 16'h8888;
    SB_DFF ootx_shift_registers_0_3_c (.Q(ootx_shift_registers_0_3), .C(clock_c), 
           .D(n11026));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i1_2_lut_3_lut_adj_740 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n217), .I3(GND_net), .O(n986));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_740.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_741 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n219), .I3(GND_net), .O(n988));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_741.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_742 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n75), .O(n972));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_742.LUT_INIT = 16'h4000;
    SB_LUT4 mod_155_add_1138_5_lut (.I0(n1610), .I1(n1610), .I2(n1631_adj_2058), 
            .I3(n22484), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1607_4 (.CI(n22609), .I0(n2311), .I1(n2324), 
            .CO(n22610));
    SB_LUT4 i1_2_lut_3_lut_adj_743 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n225), .I3(GND_net), .O(n994));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_743.LUT_INIT = 16'h4040;
    SB_DFF ootx_shift_registers_0_2_c (.Q(ootx_shift_registers_0_2), .C(clock_c), 
           .D(n11025));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 i7713_3_lut_4_lut (.I0(n942), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1223), .O(n11823));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7713_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF ootx_shift_registers_0_1_c (.Q(ootx_shift_registers_0_1), .C(clock_c), 
           .D(n11024));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_DFF ootx_shift_registers_0_0_c (.Q(ootx_shift_registers_0_0), .C(clock_c), 
           .D(n11023));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(47[9:29])
    SB_LUT4 EnabledDecoder_2_i24_2_lut_3_lut_4_lut (.I0(ootx_payloads_N_1685), 
            .I1(ootx_payloads_N_1699[0]), .I2(ootx_payloads_N_1699[1]), 
            .I3(ootx_payloads_N_1699[2]), .O(n24_adj_1903));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i24_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_adj_744 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n233), .I3(GND_net), .O(n1002));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_744.LUT_INIT = 16'h4040;
    SB_DFF i386_387_adj_745 (.Q(ootx_payloads_0_36), .C(clock_c), .D(n11022));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY counter_from_nskip_rise_640_add_4_15 (.CI(n22363), .I0(n2280), 
            .I1(counter_from_nskip_rise[13]), .CO(n22364));
    SB_DFF i284_285_adj_746 (.Q(ootx_payloads_0_2), .C(clock_c), .D(n11021));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_747 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n81), .O(n978));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_747.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_748 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n119), .O(n1016));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_748.LUT_INIT = 16'h4000;
    SB_DFF i392_393_adj_749 (.Q(ootx_payloads_0_38), .C(clock_c), .D(n11020));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_750 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n83_adj_2035), .O(n980));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_750.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_adj_751 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n249), .I3(GND_net), .O(n1018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_751.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_752 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n251), .I3(GND_net), .O(n1020));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_752.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_753 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n85), .O(n982));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_753.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_adj_754 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n255), .I3(GND_net), .O(n1024));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_754.LUT_INIT = 16'h4040;
    SB_DFFE data_484 (.Q(data), .C(clock_c), .E(n23999), .D(data_N_1765));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i1_2_lut_3_lut_adj_755 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n257), .I3(GND_net), .O(n1026));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_755.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_756 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n259), .I3(GND_net), .O(n1028));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_756.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_757 (.I0(\ootx_payloads_N_1699[8] ), .I1(\ootx_payloads_N_1699[7] ), 
            .I2(n261), .I3(GND_net), .O(n1030));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_adj_757.LUT_INIT = 16'h4040;
    SB_LUT4 mod_155_add_1875_2_lut (.I0(n2851[5]), .I1(n2851[5]), .I2(n25192), 
            .I3(VCC_net), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_355_27_lut (.I0(GND_net), .I1(\counter_from_last_rise[25] ), 
            .I2(GND_net), .I3(n22299), .O(n6340)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7121_3_lut_4_lut (.I0(n942), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_210), .O(n11231));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7121_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i365_366_adj_758 (.Q(ootx_payloads_0_29), .C(clock_c), .D(n11019));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFFESR sensor_state_switch_counter_641__i0 (.Q(sensor_state_switch_counter[0]), 
            .C(clock_c), .E(n13338), .D(n100[0]), .R(n13346));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    SB_DFF i716_717_adj_759 (.Q(ootx_payloads_0_146), .C(clock_c), .D(n11167));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_760 (.I0(n13), .I1(n24018), .I2(ootx_payloads_N_1744[1]), 
            .I3(ootx_payloads_N_1744[0]), .O(n93));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_3_lut_4_lut_adj_760.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_761 (.I0(\ootx_payloads_N_1699[8] ), 
            .I1(\ootx_payloads_N_1699[7] ), .I2(\ootx_payloads_N_1699[6] ), 
            .I3(n79), .O(n976));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i1_2_lut_3_lut_4_lut_adj_761.LUT_INIT = 16'h4000;
    SB_LUT4 i19412_2_lut_4_lut (.I0(n16_adj_2143), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24059));
    defparam i19412_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_LUT4 i19427_2_lut_4_lut (.I0(n16_adj_2143), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24089));
    defparam i19427_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 i7757_3_lut_4_lut (.I0(n1030), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1179), .O(n11867));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7757_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7165_3_lut_4_lut (.I0(n1030), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_254), .O(n11275));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7165_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7628_3_lut_4_lut (.I0(n772), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1308), .O(n11738));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7628_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i713_714_adj_762 (.Q(ootx_payloads_0_145), .C(clock_c), .D(n11166));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7036_3_lut_4_lut (.I0(n772), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_125), .O(n11146));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7036_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19411_2_lut_4_lut (.I0(n18_adj_2173), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24057));
    defparam i19411_2_lut_4_lut.LUT_INIT = 16'hce00;
    SB_DFF i710_711_adj_763 (.Q(ootx_payloads_0_144), .C(clock_c), .D(n11165));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i707_708_adj_764 (.Q(ootx_payloads_0_143), .C(clock_c), .D(n11164));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i704_705_adj_765 (.Q(ootx_payloads_0_142), .C(clock_c), .D(n11163));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i701_702_adj_766 (.Q(ootx_payloads_0_141), .C(clock_c), .D(n11162));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i698_699_adj_767 (.Q(ootx_payloads_0_140), .C(clock_c), .D(n11161));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i695_696_adj_768 (.Q(ootx_payloads_0_139), .C(clock_c), .D(n11160));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i692_693_adj_769 (.Q(ootx_payloads_0_138), .C(clock_c), .D(n11159));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i689_690_adj_770 (.Q(ootx_payloads_0_137), .C(clock_c), .D(n11158));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1607_3_lut (.I0(n2312), .I1(n2312), .I2(n2324), 
            .I3(n22608), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_3_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i287_288_adj_771 (.Q(ootx_payloads_0_3), .C(clock_c), .D(n11018));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i371_372_adj_772 (.Q(ootx_payloads_0_31), .C(clock_c), .D(n11017));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i19426_2_lut_4_lut (.I0(n18_adj_2173), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24087));
    defparam i19426_2_lut_4_lut.LUT_INIT = 16'h00ce;
    SB_LUT4 i19410_2_lut_4_lut (.I0(n19263), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24055));
    defparam i19410_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_LUT4 EnabledDecoder_2_i536_2_lut_4_lut (.I0(n88_adj_1877), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n536));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i536_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i534_2_lut_4_lut (.I0(n86_adj_1860), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n534));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i534_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_1138_5 (.CI(n22484), .I0(n1610), .I1(n1631_adj_2058), 
            .CO(n22485));
    SB_CARRY add_355_27 (.CI(n22299), .I0(\counter_from_last_rise[25] ), 
            .I1(GND_net), .CO(n22300));
    SB_LUT4 EnabledDecoder_2_i532_2_lut_4_lut (.I0(n84), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n532));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i532_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY mod_155_add_2143_9 (.CI(n22818), .I0(n3107_adj_2168), .I1(n3116), 
            .CO(n22819));
    SB_LUT4 i7712_3_lut_4_lut (.I0(n940), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1224), .O(n11822));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7712_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i663__i1 (.Q(\ootx_payload_o[0][0] ), .C(clock_c), .D(n11016));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(159[42:52])
    SB_LUT4 EnabledDecoder_2_i530_2_lut_4_lut (.I0(n82_adj_1873), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n530));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i530_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i19425_2_lut_4_lut (.I0(n19263), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24085));
    defparam i19425_2_lut_4_lut.LUT_INIT = 16'h00dc;
    SB_LUT4 EnabledDecoder_2_i528_2_lut_4_lut (.I0(n80), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n528));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i528_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i526_2_lut_4_lut (.I0(n78_adj_1891), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n526));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i526_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i524_2_lut_4_lut (.I0(n76), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n524));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i524_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF i290_291_adj_773 (.Q(ootx_payloads_0_4), .C(clock_c), .D(n11015));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 EnabledDecoder_2_i522_2_lut_4_lut (.I0(n74_adj_1899), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n522));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i522_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i67_2_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n67));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i67_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i65_2_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n65));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i65_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 EnabledDecoder_2_i114_2_lut_4_lut (.I0(n17_adj_1864), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n114_adj_2044));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i114_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i112_2_lut_4_lut (.I0(n24_adj_1903), .I1(\ootx_payloads_N_1699[3] ), 
            .I2(\ootx_payloads_N_1699[4] ), .I3(\ootx_payloads_N_1699[5] ), 
            .O(n112_adj_2043));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i112_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n63));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i63_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i19409_2_lut_4_lut (.I0(n15_adj_2148), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24053));
    defparam i19409_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_DFF i293_294_adj_774 (.Q(ootx_payloads_0_5), .C(clock_c), .D(n11014));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_15_i1_3_lut_adj_775 (.I0(payload_lengths_0_5), .I1(payload_lengths_1_5), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[5] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_15_i1_3_lut_adj_775.LUT_INIT = 16'hcaca;
    SB_LUT4 i19424_2_lut_4_lut (.I0(n15_adj_2148), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24083));
    defparam i19424_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_LUT4 Mux_14_i1_3_lut_adj_776 (.I0(payload_lengths_0_6), .I1(payload_lengths_1_6), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[6] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_14_i1_3_lut_adj_776.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_777 (.I0(n2851[16]), .I1(n1612), .I2(n1611), 
            .I3(n1610), .O(n22948));
    defparam i3_4_lut_adj_777.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_778 (.I0(n22948), .I1(n1606), .I2(n1609), .I3(GND_net), 
            .O(n16_adj_2205));
    defparam i4_3_lut_adj_778.LUT_INIT = 16'hecec;
    SB_LUT4 mod_155_add_2143_8_lut (.I0(n3108_adj_2161), .I1(n3108_adj_2161), 
            .I2(n3116), .I3(n22817), .O(n13_adj_1951)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i686_687_adj_779 (.Q(ootx_payloads_0_136), .C(clock_c), .D(n11157));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 counter_from_nskip_rise_640_add_4_14_lut (.I0(n6333[12]), .I1(n2280), 
            .I2(counter_from_nskip_rise[12]), .I3(n22362), .O(n91[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i7_4_lut_adj_780 (.I0(n1608), .I1(n1599_adj_2087), .I2(n1601_adj_2150), 
            .I3(n1598_adj_2086), .O(n19_adj_2206));
    defparam i7_4_lut_adj_780.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1875_2 (.CI(VCC_net), .I0(n2851[5]), .I1(n25192), 
            .CO(n22702));
    SB_LUT4 i7756_3_lut_4_lut (.I0(n1028), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1180), .O(n11866));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7756_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i683_684_adj_781 (.Q(ootx_payloads_0_135), .C(clock_c), .D(n11156));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i6_2_lut_adj_782 (.I0(n1607), .I1(n1602_adj_2154), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_2207));
    defparam i6_2_lut_adj_782.LUT_INIT = 16'heeee;
    SB_LUT4 i7164_3_lut_4_lut (.I0(n1028), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_253), .O(n11274));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7164_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_783 (.I0(n19_adj_2206), .I1(n1604), .I2(n16_adj_2205), 
            .I3(n1600_adj_2090), .O(n22_adj_2208));
    defparam i10_4_lut_adj_783.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_7_Mux_1_i1_3_lut (.I0(\ootx_states[0] [1]), .I1(\ootx_states[1] [1]), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1744[1]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[21:31])
    defparam mux_7_Mux_1_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i680_681_adj_784 (.Q(ootx_payloads_0_134), .C(clock_c), .D(n11155));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1138_4_lut (.I0(n1611), .I1(n1611), .I2(n1631_adj_2058), 
            .I3(n22483), .O(n1710)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_785 (.I0(n1603), .I1(n22_adj_2208), .I2(n18_adj_2207), 
            .I3(n1605), .O(n1631_adj_2058));
    defparam i11_4_lut_adj_785.LUT_INIT = 16'hfffe;
    SB_DFF i677_678_adj_786 (.Q(ootx_payloads_0_133), .C(clock_c), .D(n11154));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_13_i1_3_lut_adj_787 (.I0(payload_lengths_0_7), .I1(payload_lengths_1_7), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[7] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_13_i1_3_lut_adj_787.LUT_INIT = 16'hcaca;
    SB_LUT4 i7627_3_lut_4_lut (.I0(n770), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1309), .O(n11737));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7627_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i368_369_adj_788 (.Q(ootx_payloads_0_30), .C(clock_c), .D(n11013));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_12_i1_3_lut_adj_789 (.I0(payload_lengths_0_8), .I1(payload_lengths_1_8), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[8] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_12_i1_3_lut_adj_789.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_11_i1_3_lut_adj_790 (.I0(payload_lengths_0_9), .I1(payload_lengths_1_9), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[9] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_11_i1_3_lut_adj_790.LUT_INIT = 16'hcaca;
    SB_LUT4 i7035_3_lut_4_lut (.I0(n770), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_124), .O(n11145));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7035_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_7_Mux_0_i1_3_lut (.I0(\ootx_states[0] [0]), .I1(\ootx_states[1][0] ), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(ootx_payloads_N_1744[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(86[21:31])
    defparam mux_7_Mux_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7120_3_lut_4_lut (.I0(n940), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_209), .O(n11230));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7120_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_14 (.CI(n22362), .I0(n2280), 
            .I1(counter_from_nskip_rise[12]), .CO(n22363));
    SB_CARRY mod_155_add_1607_3 (.CI(n22608), .I0(n2312), .I1(n2324), 
            .CO(n22609));
    SB_LUT4 i19408_2_lut_4_lut (.I0(n17_adj_2144), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24051));
    defparam i19408_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i20529_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25197));
    defparam i20529_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_155_add_1607_2_lut (.I0(n2851[9]), .I1(n2851[9]), .I2(n25198), 
            .I3(VCC_net), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFF ootx_crc32_2_o_i0_i0 (.Q(\ootx_crc32_o[1] [0]), .C(clock_c), 
           .D(n11012));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 Mux_10_i1_3_lut_adj_791 (.I0(payload_lengths_0_10), .I1(payload_lengths_1_10), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[10] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_10_i1_3_lut_adj_791.LUT_INIT = 16'hcaca;
    SB_DFF ootx_crc32_1_o_i0_i0 (.Q(\ootx_crc32_o[0] [0]), .C(clock_c), 
           .D(n11011));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 Mux_9_i1_3_lut_adj_792 (.I0(payload_lengths_0_11), .I1(payload_lengths_1_11), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(\ootx_payloads_N_1730[11] ));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_9_i1_3_lut_adj_792.LUT_INIT = 16'hcaca;
    SB_LUT4 i19423_2_lut_4_lut (.I0(n17_adj_2144), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24081));
    defparam i19423_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_DFF i296_297_adj_793 (.Q(ootx_payloads_0_6), .C(clock_c), .D(n11010));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i2_2_lut_adj_794 (.I0(n2312), .I1(n2310), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_2209));
    defparam i2_2_lut_adj_794.LUT_INIT = 16'heeee;
    SB_LUT4 i15211_4_lut (.I0(n2851[9]), .I1(n2309), .I2(n6_adj_2209), 
            .I3(n2311), .O(n19307));
    defparam i15211_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i11_4_lut_adj_795 (.I0(n2299), .I1(n2296), .I2(n19307), .I3(n2293), 
            .O(n30_adj_2210));
    defparam i11_4_lut_adj_795.LUT_INIT = 16'hfffe;
    SB_DFF i362_363_adj_796 (.Q(ootx_payloads_0_28), .C(clock_c), .D(n11009));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i15_4_lut_adj_797 (.I0(n2295), .I1(n30_adj_2210), .I2(n2298), 
            .I3(n2305), .O(n34_adj_2211));
    defparam i15_4_lut_adj_797.LUT_INIT = 16'hfffe;
    SB_DFF i299_300_adj_798 (.Q(ootx_payloads_0_7), .C(clock_c), .D(n11008));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i13_4_lut_adj_799 (.I0(n2300), .I1(n2292), .I2(n2302), .I3(n2291), 
            .O(n32_adj_2212));
    defparam i13_4_lut_adj_799.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_800 (.I0(n2307), .I1(n2308), .I2(n2301), .I3(n2294), 
            .O(n33_adj_2213));
    defparam i14_4_lut_adj_800.LUT_INIT = 16'hfffe;
    SB_DFFR ootx_states_0__i0_i0 (.Q(\ootx_states[0] [0]), .C(clock_c), 
            .D(n25), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i12_4_lut_adj_801 (.I0(n2303), .I1(n2306), .I2(n2304), .I3(n2297), 
            .O(n31_adj_2215));
    defparam i12_4_lut_adj_801.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_802 (.I0(n31_adj_2215), .I1(n33_adj_2213), .I2(n32_adj_2212), 
            .I3(n34_adj_2211), .O(n2324));
    defparam i18_4_lut_adj_802.LUT_INIT = 16'hfffe;
    SB_LUT4 EnabledDecoder_2_i61_2_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n61));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i61_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFF i302_303_adj_803 (.Q(ootx_payloads_0_8), .C(clock_c), .D(n11006));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i19407_2_lut_4_lut (.I0(n19_adj_2172), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24049));
    defparam i19407_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i19422_2_lut_4_lut (.I0(n19_adj_2172), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24079));
    defparam i19422_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_CARRY mod_155_add_1138_4 (.CI(n22483), .I0(n1611), .I1(n1631_adj_2058), 
            .CO(n22484));
    SB_LUT4 i7755_3_lut_4_lut (.I0(n1026), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1181), .O(n11865));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7755_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_355_26_lut (.I0(GND_net), .I1(\counter_from_last_rise[24] ), 
            .I2(GND_net), .I3(n22298), .O(n6341)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7163_3_lut_4_lut (.I0(n1026), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_252), .O(n11273));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7163_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i305_306_adj_804 (.Q(ootx_payloads_0_9), .C(clock_c), .D(n11005));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 EnabledDecoder_2_i258_2_lut_3_lut (.I0(n65_c), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n258));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i258_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 counter_from_nskip_rise_640_add_4_13_lut (.I0(n6333[11]), .I1(n2280), 
            .I2(counter_from_nskip_rise[11]), .I3(n22361), .O(n91[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 EnabledDecoder_2_i257_2_lut_3_lut (.I0(n65_c), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n257));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i257_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7754_3_lut_4_lut (.I0(n1024), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1182), .O(n11864));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7754_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7162_3_lut_4_lut (.I0(n1024), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_251), .O(n11272));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7162_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i308_309_adj_805 (.Q(ootx_payloads_0_10), .C(clock_c), .D(n11004));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i19406_2_lut_4_lut (.I0(n12_adj_2180), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24047));
    defparam i19406_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i19421_2_lut_4_lut (.I0(n12_adj_2180), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24077));
    defparam i19421_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_DFF i311_312_adj_806 (.Q(ootx_payloads_0_11), .C(clock_c), .D(n11003));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7753_3_lut_4_lut (.I0(n1022), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1183), .O(n11863));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7753_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 ootx_payloads_I_14_i3_2_lut (.I0(ootx_payloads_N_1744[0]), .I1(ootx_payloads_N_1744[1]), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(140[13:44])
    defparam ootx_payloads_I_14_i3_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n59));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i59_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i7161_3_lut_4_lut (.I0(n1022), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_250), .O(n11271));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7161_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_807 (.I0(n93), .I1(new_data), .I2(reset_c), 
            .I3(GND_net), .O(n20123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_3_lut_adj_807.LUT_INIT = 16'h0808;
    SB_LUT4 i7752_3_lut_4_lut (.I0(n1020), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1184), .O(n11862));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7752_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i57_2_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n57));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i57_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i7160_3_lut_4_lut (.I0(n1020), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_249), .O(n11270));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7160_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i55_2_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n55));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i55_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY mod_155_add_2076_5 (.CI(n22785), .I0(n3010), .I1(n3017), 
            .CO(n22786));
    SB_LUT4 mod_155_add_1138_3_lut (.I0(n1612), .I1(n1612), .I2(n1631_adj_2058), 
            .I3(n22482), .O(n1711)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_3_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_26 (.CI(n22298), .I0(\counter_from_last_rise[24] ), 
            .I1(GND_net), .CO(n22299));
    SB_LUT4 mod_155_add_2076_4_lut (.I0(n3011), .I1(n3011), .I2(n3017), 
            .I3(n22784), .O(n3110_adj_2159)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2143_8 (.CI(n22817), .I0(n3108_adj_2161), .I1(n3116), 
            .CO(n22818));
    SB_CARRY counter_from_nskip_rise_640_add_4_13 (.CI(n22361), .I0(n2280), 
            .I1(counter_from_nskip_rise[11]), .CO(n22362));
    SB_LUT4 EnabledDecoder_2_i53_2_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n53));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i53_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY mod_155_add_1607_2 (.CI(VCC_net), .I0(n2851[9]), .I1(n25198), 
            .CO(n22608));
    SB_DFF i674_675_adj_808 (.Q(ootx_payloads_0_132), .C(clock_c), .D(n11153));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i19405_2_lut_4_lut (.I0(n14_adj_2149), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24045));
    defparam i19405_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i19420_2_lut_4_lut (.I0(n14_adj_2149), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24075));
    defparam i19420_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_LUT4 i7008_3_lut_4_lut (.I0(n716), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_97), .O(n11118));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7008_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7600_3_lut_4_lut (.I0(n716), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1336), .O(n11710));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7600_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7751_3_lut_4_lut (.I0(n1018), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1185), .O(n11861));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7751_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i671_672_adj_809 (.Q(ootx_payloads_0_131), .C(clock_c), .D(n11152));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7159_3_lut_4_lut (.I0(n1018), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_248), .O(n11269));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7159_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6948_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_16), .I3(ootx_shift_registers_1_17), 
            .O(n11058));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6948_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i314_315_adj_810 (.Q(ootx_payloads_0_12), .C(clock_c), .D(n11002));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_2143_7_lut (.I0(n3109_adj_2162), .I1(n3109_adj_2162), 
            .I2(n25181), .I3(n22816), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_7_lut.LUT_INIT = 16'hA3AC;
    SB_DFF i317_318_adj_811 (.Q(ootx_payloads_0_13), .C(clock_c), .D(n11001));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1942_26 (.CI(n22751), .I0(n2789), .I1(n2819), 
            .CO(n22752));
    SB_LUT4 i1_4_lut_4_lut (.I0(reset_c), .I1(sensor_state_switch_counter[0]), 
            .I2(n10_adj_2057), .I3(sensor_state_switch_counter[4]), .O(n13338));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5554;
    SB_DFF i377_378_adj_812 (.Q(ootx_payloads_0_33), .C(clock_c), .D(n11000));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1808_27_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n22701), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_7_i1_3_lut_adj_813 (.I0(payload_lengths_0_13), .I1(payload_lengths_1_13), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n577[13]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_7_i1_3_lut_adj_813.LUT_INIT = 16'hcaca;
    SB_LUT4 add_355_25_lut (.I0(GND_net), .I1(\counter_from_last_rise[23] ), 
            .I2(GND_net), .I3(n22297), .O(n6342)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_155_add_1540_23_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n22607), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15169_2_lut_4_lut (.I0(ootx_payloads_N_1699[0]), .I1(n88), 
            .I2(ootx_payloads_N_1699[1]), .I3(ootx_payloads_N_1699[2]), 
            .O(n19263));
    defparam i15169_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 EnabledDecoder_2_i535_2_lut_4_lut (.I0(n88_adj_1877), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n535));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i535_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 EnabledDecoder_2_i68_2_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n68));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i68_2_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i533_2_lut_4_lut (.I0(n86_adj_1860), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n533));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i533_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 EnabledDecoder_2_i66_2_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n66));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i66_2_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i64_2_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n64));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i64_2_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i62_2_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n62));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i62_2_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i60_2_lut_4_lut (.I0(n11_adj_2070), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n60));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i60_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i531_2_lut_4_lut (.I0(n84), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n531));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i531_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_CARRY mod_155_add_1138_3 (.CI(n22482), .I0(n1612), .I1(n1631_adj_2058), 
            .CO(n22483));
    SB_CARRY mod_155_add_2076_4 (.CI(n22784), .I0(n3011), .I1(n3017), 
            .CO(n22785));
    SB_LUT4 mod_155_add_1942_25_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n22750), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 EnabledDecoder_2_i58_2_lut_4_lut (.I0(n9), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n58));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i58_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 counter_from_nskip_rise_640_add_4_12_lut (.I0(n6355), .I1(n2280), 
            .I2(counter_from_nskip_rise[10]), .I3(n22360), .O(n91[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_355_25 (.CI(n22297), .I0(\counter_from_last_rise[23] ), 
            .I1(GND_net), .CO(n22298));
    SB_LUT4 EnabledDecoder_2_i56_2_lut_4_lut (.I0(n12_adj_2072), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n56));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i56_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i54_2_lut_4_lut (.I0(n10_adj_2079), .I1(ootx_payloads_N_1699[2]), 
            .I2(\ootx_payloads_N_1699[3] ), .I3(\ootx_payloads_N_1699[4] ), 
            .O(n54));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(173[29:54])
    defparam EnabledDecoder_2_i54_2_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i529_2_lut_4_lut (.I0(n82_adj_1873), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n529));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i529_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mod_155_add_1138_2_lut (.I0(n2851[16]), .I1(n2851[16]), .I2(n25199), 
            .I3(VCC_net), .O(n1712)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 EnabledDecoder_2_i527_2_lut_4_lut (.I0(n80), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n527));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i527_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_CARRY mod_155_add_1942_25 (.CI(n22750), .I0(n2790), .I1(n2819), 
            .CO(n22751));
    SB_LUT4 EnabledDecoder_2_i525_2_lut_4_lut (.I0(n78_adj_1891), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n525));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i525_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 EnabledDecoder_2_i523_2_lut_4_lut (.I0(n76), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n523));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i523_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mod_155_add_2076_3_lut (.I0(n3012), .I1(n3012), .I2(n3017), 
            .I3(n22783), .O(n3111_adj_2158)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_3_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 Mux_6_i1_3_lut_adj_814 (.I0(payload_lengths_0_14), .I1(payload_lengths_1_14), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n577[14]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_6_i1_3_lut_adj_814.LUT_INIT = 16'hcaca;
    SB_CARRY counter_from_nskip_rise_640_add_4_12 (.CI(n22360), .I0(n2280), 
            .I1(counter_from_nskip_rise[10]), .CO(n22361));
    SB_LUT4 EnabledDecoder_2_i20_2_lut_3_lut_4_lut (.I0(ootx_payloads_N_1685), 
            .I1(ootx_payloads_N_1699[0]), .I2(ootx_payloads_N_1699[1]), 
            .I3(ootx_payloads_N_1699[2]), .O(n20_adj_1943));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i20_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 mod_155_add_1808_26_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n22700), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6932_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_0), .I3(ootx_shift_registers_1_1), 
            .O(n11042));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6932_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n13329), .I1(reset_c), .I2(sensor_N_132), 
            .I3(sensor_state), .O(n23693));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hdf02;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_4_lut (.I0(ootx_payloads_N_1699[0]), 
            .I1(n88), .I2(ootx_payloads_N_1699[1]), .I3(ootx_payloads_N_1699[2]), 
            .O(n12_adj_2180));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(119[37:62])
    defparam EnabledDecoder_2_i12_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFF i668_669_adj_815 (.Q(ootx_payloads_0_130), .C(clock_c), .D(n11151));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_816 (.I0(n13329), .I1(reset_c), .I2(sensor_N_132), 
            .I3(sensor_state), .O(n13346));
    defparam i1_2_lut_3_lut_4_lut_adj_816.LUT_INIT = 16'h2002;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(n13329), .I1(reset_c), .I2(sensor_N_132), 
            .I3(n23997), .O(n23999));
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i521_2_lut_4_lut (.I0(n74_adj_1899), .I1(\ootx_payloads_N_1699[6] ), 
            .I2(\ootx_payloads_N_1699[7] ), .I3(\ootx_payloads_N_1699[8] ), 
            .O(n521));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i521_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_CARRY mod_155_add_2143_7 (.CI(n22816), .I0(n3109_adj_2162), .I1(n25181), 
            .CO(n22817));
    SB_LUT4 PrioSelect_81_i2_3_lut_4_lut (.I0(data), .I1(n4501), .I2(n432), 
            .I3(\lighthouse[0] ), .O(n114));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_81_i2_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 mod_155_add_1540_22_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n22606), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1540_22 (.CI(n22606), .I0(n2193), .I1(n2225), 
            .CO(n22607));
    SB_LUT4 i1_3_lut_4_lut_adj_817 (.I0(counter_from_nskip_rise[1]), .I1(counter_from_nskip_rise[4]), 
            .I2(counter_from_nskip_rise[2]), .I3(counter_from_nskip_rise[3]), 
            .O(n6_adj_1934));
    defparam i1_3_lut_4_lut_adj_817.LUT_INIT = 16'hccc8;
    SB_LUT4 i3_2_lut_adj_818 (.I0(n2502), .I1(n2501), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_2226));
    defparam i3_2_lut_adj_818.LUT_INIT = 16'heeee;
    SB_CARRY mod_155_add_1138_2 (.CI(VCC_net), .I0(n2851[16]), .I1(n25199), 
            .CO(n22482));
    SB_LUT4 i2_3_lut_4_lut_adj_819 (.I0(counter_from_last_rise[2]), .I1(counter_from_last_rise_c[5]), 
            .I2(counter_from_last_rise[4]), .I3(counter_from_last_rise[3]), 
            .O(n22900));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(40[9:31])
    defparam i2_3_lut_4_lut_adj_819.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_820 (.I0(n2494), .I1(n2503), .I2(n2497), .I3(n2491), 
            .O(n34_adj_2227));
    defparam i13_4_lut_adj_820.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_821 (.I0(\lighthouse[0] ), .I1(n93), .I2(n23989), 
            .I3(n4729), .O(n23991));
    defparam i1_3_lut_4_lut_adj_821.LUT_INIT = 16'hf080;
    SB_LUT4 i11_3_lut_adj_822 (.I0(n2506), .I1(n2492), .I2(n2489), .I3(GND_net), 
            .O(n32_adj_2228));
    defparam i11_3_lut_adj_822.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_823 (.I0(n2851[7]), .I1(n2512), .I2(n2511), .I3(n2510), 
            .O(n22895));
    defparam i3_4_lut_adj_823.LUT_INIT = 16'hfffe;
    SB_LUT4 counter_from_nskip_rise_640_add_4_11_lut (.I0(n6356), .I1(n2280), 
            .I2(counter_from_nskip_rise[9]), .I3(n22359), .O(n91[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_355_24_lut (.I0(GND_net), .I1(\counter_from_last_rise[22] ), 
            .I2(GND_net), .I3(n22296), .O(n6343)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_824 (.I0(new_data), .I1(reset_c), .I2(n24110), 
            .I3(GND_net), .O(n1119));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i1_2_lut_3_lut_adj_824.LUT_INIT = 16'h0202;
    SB_LUT4 i17_4_lut_adj_825 (.I0(n2490), .I1(n34_adj_2227), .I2(n24_adj_2226), 
            .I3(n2508), .O(n38_adj_2229));
    defparam i17_4_lut_adj_825.LUT_INIT = 16'hfffe;
    SB_DFF i665_666_adj_826 (.Q(ootx_payloads_0_129), .C(clock_c), .D(n11150));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i19444_2_lut_4_lut (.I0(ootx_payloads_N_1744[0]), .I1(ootx_payloads_N_1744[1]), 
            .I2(n2679), .I3(n2680), .O(n24110));
    defparam i19444_2_lut_4_lut.LUT_INIT = 16'hbbfb;
    SB_LUT4 i15_4_lut_adj_827 (.I0(n2500), .I1(n2505), .I2(n2496), .I3(n2493), 
            .O(n36_adj_2230));
    defparam i15_4_lut_adj_827.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_155_add_1071_16_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n22481), .O(n1598_adj_2086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_16_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i320_321_adj_828 (.Q(ootx_payloads_0_14), .C(clock_c), .D(n10999));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i16_4_lut_adj_829 (.I0(n22895), .I1(n32_adj_2228), .I2(n2504), 
            .I3(n2509), .O(n37_adj_2231));
    defparam i16_4_lut_adj_829.LUT_INIT = 16'hfefc;
    SB_DFF i662_663_adj_830 (.Q(ootx_payloads_0_128), .C(clock_c), .D(n11149));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i14803_2_lut_3_lut (.I0(n35), .I1(reset_c), .I2(n4729), .I3(GND_net), 
            .O(data_counters_N_1776));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i14803_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFF i659_660_adj_831 (.Q(ootx_payloads_0_127), .C(clock_c), .D(n11148));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i323_324_adj_832 (.Q(ootx_payloads_0_15), .C(clock_c), .D(n10998));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 Mux_5_i1_3_lut (.I0(payload_lengths_0_15), .I1(payload_lengths_1_15), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n577[15]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(142[66:76])
    defparam Mux_5_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i864_2_lut (.I0(sensor_N_132), .I1(sensor_state), .I2(GND_net), 
            .I3(GND_net), .O(n2276));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(199[5] 341[12])
    defparam i864_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6947_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_15), .I3(ootx_shift_registers_1_16), 
            .O(n11057));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6947_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i656_657_adj_833 (.Q(ootx_payloads_0_126), .C(clock_c), .D(n11147));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i653_654_adj_834 (.Q(ootx_payloads_0_125), .C(clock_c), .D(n11146));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i14_4_lut_adj_835 (.I0(n2498), .I1(n2495), .I2(n2507), .I3(n2499), 
            .O(n35_adj_2232));
    defparam i14_4_lut_adj_835.LUT_INIT = 16'hfffe;
    SB_LUT4 PrioSelect_145_i2_3_lut_4_lut (.I0(data), .I1(n4501), .I2(n432), 
            .I3(\lighthouse[0] ), .O(n178));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(58[9:24])
    defparam PrioSelect_145_i2_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY counter_from_nskip_rise_640_add_4_11 (.CI(n22359), .I0(n2280), 
            .I1(counter_from_nskip_rise[9]), .CO(n22360));
    SB_LUT4 i20336_2_lut_3_lut (.I0(n13329), .I1(sensor_N_132), .I2(sensor_state), 
            .I3(GND_net), .O(n24697));
    defparam i20336_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_CARRY add_355_24 (.CI(n22296), .I0(\counter_from_last_rise[22] ), 
            .I1(GND_net), .CO(n22297));
    SB_LUT4 i20185_2_lut_4_lut (.I0(n2679), .I1(n2680), .I2(data), .I3(n13), 
            .O(n24564));
    defparam i20185_2_lut_4_lut.LUT_INIT = 16'hdfdd;
    SB_LUT4 i20_4_lut_adj_836 (.I0(n35_adj_2232), .I1(n37_adj_2231), .I2(n36_adj_2230), 
            .I3(n38_adj_2229), .O(n2522));
    defparam i20_4_lut_adj_836.LUT_INIT = 16'hfffe;
    SB_LUT4 i19404_2_lut_4_lut (.I0(n16_adj_2143), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24043));
    defparam i19404_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_DFF i326_327_adj_837 (.Q(ootx_payloads_0_16), .C(clock_c), .D(n10997));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1808_26 (.CI(n22700), .I0(n2589), .I1(n2621), 
            .CO(n22701));
    SB_LUT4 i19419_2_lut_4_lut (.I0(n16_adj_2143), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24073));
    defparam i19419_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_LUT4 mod_155_add_1540_21_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n22605), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7750_3_lut_4_lut (.I0(n1016), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1186), .O(n11860));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7750_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7158_3_lut_4_lut (.I0(n1016), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_247), .O(n11268));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7158_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19403_2_lut_4_lut (.I0(n18_adj_2173), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24041));
    defparam i19403_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_adj_838 (.I0(n22943), .I1(n9513), .I2(GND_net), .I3(GND_net), 
            .O(n2283));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(69[3] 344[10])
    defparam i1_2_lut_adj_838.LUT_INIT = 16'h4444;
    SB_LUT4 i5_3_lut_adj_839 (.I0(n1306_c), .I1(n1307_c), .I2(n1303_c), 
            .I3(GND_net), .O(n14_adj_2233));
    defparam i5_3_lut_adj_839.LUT_INIT = 16'hfefe;
    SB_LUT4 i6946_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_14), .I3(ootx_shift_registers_1_15), 
            .O(n11056));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6946_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i19418_2_lut_4_lut (.I0(n18_adj_2173), .I1(n432), .I2(\ootx_payloads_N_1699[3] ), 
            .I3(\lighthouse[0] ), .O(n24071));
    defparam i19418_2_lut_4_lut.LUT_INIT = 16'h00ec;
    SB_CARRY mod_155_add_1540_21 (.CI(n22605), .I0(n2194), .I1(n2225), 
            .CO(n22606));
    SB_LUT4 i20487_3_lut_4_lut (.I0(ootx_payloads_N_1744[1]), .I1(ootx_payloads_N_1744[0]), 
            .I2(n35), .I3(new_data), .O(n4731));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i20487_3_lut_4_lut.LUT_INIT = 16'h01ff;
    SB_LUT4 i3_4_lut_adj_840 (.I0(n2851[19]), .I1(n1312_adj_1925), .I2(n1311_adj_1923), 
            .I3(n1310_c), .O(n22872));
    defparam i3_4_lut_adj_840.LUT_INIT = 16'hfffe;
    SB_LUT4 i6945_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_13), .I3(ootx_shift_registers_1_14), 
            .O(n11055));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6945_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_841 (.I0(ootx_payloads_N_1744[1]), .I1(ootx_payloads_N_1744[0]), 
            .I2(new_data), .I3(GND_net), .O(n9989));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    defparam i1_2_lut_3_lut_adj_841.LUT_INIT = 16'hefef;
    SB_LUT4 i3_2_lut_adj_842 (.I0(n1305_c), .I1(n1304_c), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_2234));
    defparam i3_2_lut_adj_842.LUT_INIT = 16'heeee;
    SB_DFF i329_330_adj_843 (.Q(ootx_payloads_0_17), .C(clock_c), .D(n10996));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7749_3_lut_4_lut (.I0(n1014), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1187), .O(n11859));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7749_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7157_3_lut_4_lut (.I0(n1014), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_246), .O(n11267));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7157_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i20197_2_lut_3_lut (.I0(\counter_from_last_rise[8] ), .I1(counter_from_last_rise[2]), 
            .I2(counter_from_last_rise[3]), .I3(GND_net), .O(n24682));
    defparam i20197_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_844 (.I0(ootx_payloads_N_1744[1]), .I1(data), 
            .I2(n13), .I3(n30), .O(n31));
    defparam i1_3_lut_4_lut_adj_844.LUT_INIT = 16'h20aa;
    SB_LUT4 i7_4_lut_adj_845 (.I0(n22872), .I1(n14_adj_2233), .I2(n1301_c), 
            .I3(n1309_c), .O(n16_adj_2235));
    defparam i7_4_lut_adj_845.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_155_add_1071_15_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n22480), .O(n1599_adj_2087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i395_396_adj_846 (.Q(ootx_payloads_0_39), .C(clock_c), .D(n10995));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 add_355_23_lut (.I0(GND_net), .I1(\counter_from_last_rise[21] ), 
            .I2(GND_net), .I3(n22295), .O(n6344)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut_adj_847 (.I0(n1308_c), .I1(n16_adj_2235), .I2(n12_adj_2234), 
            .I3(n1302_c), .O(n1334_c));
    defparam i8_4_lut_adj_847.LUT_INIT = 16'hfffe;
    SB_LUT4 i20305_2_lut_3_lut (.I0(\counter_from_last_rise[8] ), .I1(counter_from_last_rise[2]), 
            .I2(counter_from_last_rise[1]), .I3(GND_net), .O(n24674));
    defparam i20305_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_848 (.I0(\counter_from_last_rise[8] ), .I1(\counter_from_last_rise[6] ), 
            .I2(\counter_from_last_rise[7] ), .I3(GND_net), .O(n4_adj_1917));
    defparam i1_2_lut_3_lut_adj_848.LUT_INIT = 16'h8080;
    SB_LUT4 Mux_33_i1_3_lut_adj_849 (.I0(bit_counters_0_3), .I1(bit_counters_1_3), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[3]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_33_i1_3_lut_adj_849.LUT_INIT = 16'hcaca;
    SB_LUT4 Mux_32_i1_3_lut_adj_850 (.I0(bit_counters_0_4), .I1(bit_counters_1_4), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[4]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_32_i1_3_lut_adj_850.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_from_nskip_rise_640_add_4_10_lut (.I0(n6357), .I1(n2280), 
            .I2(counter_from_nskip_rise[8]), .I3(n22358), .O(n91[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mod_155_add_1071_15 (.CI(n22480), .I0(n1500), .I1(n1532), 
            .CO(n22481));
    SB_LUT4 Mux_275_i1_3_lut (.I0(ootx_payloads_0_0), .I1(ootx_payloads_1_0), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2[0]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(162[42:52])
    defparam Mux_275_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13560_4_lut_4_lut (.I0(\counter_from_last_rise[8] ), .I1(\counter_from_last_rise[6] ), 
            .I2(\counter_from_last_rise[7] ), .I3(n24676), .O(n223));
    defparam i13560_4_lut_4_lut.LUT_INIT = 16'ha8a0;
    SB_DFF i332_333_adj_851 (.Q(ootx_payloads_0_18), .C(clock_c), .D(n10994));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i13601_3_lut_4_lut (.I0(\counter_from_last_rise[8] ), .I1(\counter_from_last_rise[6] ), 
            .I2(counter_from_last_rise_c[5]), .I3(n119_adj_2050), .O(n193_adj_2051));
    defparam i13601_3_lut_4_lut.LUT_INIT = 16'hf808;
    SB_CARRY counter_from_nskip_rise_640_add_4_10 (.CI(n22358), .I0(n2280), 
            .I1(counter_from_nskip_rise[8]), .CO(n22359));
    SB_CARRY add_355_23 (.CI(n22295), .I0(\counter_from_last_rise[21] ), 
            .I1(GND_net), .CO(n22296));
    SB_LUT4 i7748_3_lut_4_lut (.I0(n1012), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1188), .O(n11858));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7748_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i335_336_adj_852 (.Q(ootx_payloads_0_19), .C(clock_c), .D(n10993));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1808_25_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n22699), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_25_lut.LUT_INIT = 16'hCA3A;
    SB_DFF i338_339_adj_853 (.Q(ootx_payloads_0_20), .C(clock_c), .D(n10992));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7156_3_lut_4_lut (.I0(n1012), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_245), .O(n11266));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7156_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7747_3_lut_4_lut (.I0(n1010), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1189), .O(n11857));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7747_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7155_3_lut_4_lut (.I0(n1010), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_244), .O(n11265));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7155_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i341_342_adj_854 (.Q(ootx_payloads_0_21), .C(clock_c), .D(n10991));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1540_20_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n22604), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1808_25 (.CI(n22699), .I0(n2590), .I1(n2621), 
            .CO(n22700));
    SB_LUT4 i20510_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25178));
    defparam i20510_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7746_3_lut_4_lut (.I0(n1008), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1190), .O(n11856));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7746_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i374_375_adj_855 (.Q(ootx_payloads_0_32), .C(clock_c), .D(n10990));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i20516_1_lut (.I0(n1433_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25184));
    defparam i20516_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7154_3_lut_4_lut (.I0(n1008), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_243), .O(n11264));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7154_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2143_6_lut (.I0(n3110_adj_2159), .I1(n3110_adj_2159), 
            .I2(n3116), .I3(n22815), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_155_add_1071_14_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n22479), .O(n1600_adj_2090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1540_20 (.CI(n22604), .I0(n2195), .I1(n2225), 
            .CO(n22605));
    SB_LUT4 i7017_3_lut_4_lut (.I0(n734), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_106), .O(n11127));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7017_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7609_3_lut_4_lut (.I0(n734), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1327), .O(n11719));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7609_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i344_345_adj_856 (.Q(ootx_payloads_0_22), .C(clock_c), .D(n10989));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_DFF i347_348_adj_857 (.Q(ootx_payloads_0_23), .C(clock_c), .D(n10988));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i6992_3_lut_4_lut (.I0(n684), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_81), .O(n11102));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6972_3_lut_4_lut (.I0(n644), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_61), .O(n11082));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6972_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 counter_from_nskip_rise_640_add_4_9_lut (.I0(n6358), .I1(n2280), 
            .I2(counter_from_nskip_rise[7]), .I3(n22357), .O(n91[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_9_lut.LUT_INIT = 16'h8BB8;
    SB_DFF i350_351_adj_858 (.Q(ootx_payloads_0_24), .C(clock_c), .D(n10987));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_1071_14 (.CI(n22479), .I0(n1501), .I1(n1532), 
            .CO(n22480));
    SB_LUT4 i7707_3_lut_4_lut (.I0(n930), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1229), .O(n11817));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7707_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_355_22_lut (.I0(GND_net), .I1(\counter_from_last_rise[20] ), 
            .I2(GND_net), .I3(n22294), .O(n6345)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7584_3_lut_4_lut (.I0(n684), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1352), .O(n11694));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7584_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFR ootx_states_1__i0_i0 (.Q(\ootx_states[1][0] ), .C(clock_c), 
            .D(n20_adj_33), .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut (.I0(n29_adj_1852), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n94_adj_1872));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i94_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_CARRY mod_155_add_2143_6 (.CI(n22815), .I0(n3110_adj_2159), .I1(n3116), 
            .CO(n22816));
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut (.I0(n29_adj_1852), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n93_adj_2014));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i93_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i7016_3_lut_4_lut (.I0(n732), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_105), .O(n11126));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7016_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY counter_from_nskip_rise_640_add_4_9 (.CI(n22357), .I0(n2280), 
            .I1(counter_from_nskip_rise[7]), .CO(n22358));
    SB_LUT4 i10_4_lut_adj_859 (.I0(n2204), .I1(n2198), .I2(n2194), .I3(n2207), 
            .O(n28_adj_2237));
    defparam i10_4_lut_adj_859.LUT_INIT = 16'hfffe;
    SB_CARRY add_355_22 (.CI(n22294), .I0(\counter_from_last_rise[20] ), 
            .I1(GND_net), .CO(n22295));
    SB_LUT4 i7608_3_lut_4_lut (.I0(n732), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1328), .O(n11718));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7608_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i220_2_lut_3_lut (.I0(n60_adj_2038), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n220));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i220_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i380_381_adj_860 (.Q(ootx_payloads_0_34), .C(clock_c), .D(n10985));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_2143_5_lut (.I0(n3111_adj_2158), .I1(n3111_adj_2158), 
            .I2(n3116), .I3(n22814), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2076_3 (.CI(n22783), .I0(n3012), .I1(n3017), 
            .CO(n22784));
    SB_LUT4 mod_155_add_1540_19_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n22603), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6944_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_12), .I3(ootx_shift_registers_1_13), 
            .O(n11054));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6944_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i219_2_lut_3_lut (.I0(n60_adj_2038), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n219));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i219_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i172_2_lut_3_lut (.I0(n43_adj_1944), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n172));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i172_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i171_2_lut_3_lut (.I0(n43_adj_1944), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n171));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i171_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i7745_3_lut_4_lut (.I0(n1006), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1191), .O(n11855));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7745_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i353_354_adj_861 (.Q(ootx_payloads_0_25), .C(clock_c), .D(n10984));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2143_5 (.CI(n22814), .I0(n3111_adj_2158), .I1(n3116), 
            .CO(n22815));
    SB_LUT4 EnabledDecoder_2_i90_2_lut (.I0(n58_adj_2048), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n90_adj_1876));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i90_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7153_3_lut_4_lut (.I0(n1006), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_242), .O(n11263));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7153_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mod_155_add_2076_2_lut (.I0(n2851[2]), .I1(n2851[2]), .I2(n25183), 
            .I3(VCC_net), .O(n3112_c)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_355_21_lut (.I0(GND_net), .I1(\counter_from_last_rise[19] ), 
            .I2(GND_net), .I3(n22293), .O(n6346)) /* synthesis syn_instantiated=1 */ ;
    defparam add_355_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7115_3_lut_4_lut (.I0(n930), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_204), .O(n11225));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7115_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7015_3_lut_4_lut (.I0(n730), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_104), .O(n11125));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7015_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7607_3_lut_4_lut (.I0(n730), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1329), .O(n11717));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7607_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i356_357_adj_862 (.Q(ootx_payloads_0_26), .C(clock_c), .D(n10983));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 EnabledDecoder_2_i218_2_lut_3_lut (.I0(n58_adj_2048), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n218));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i218_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i217_2_lut_3_lut (.I0(n58_adj_2048), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n217));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i217_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7744_3_lut_4_lut (.I0(n1004), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1192), .O(n11854));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7744_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i20526_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n25194));
    defparam i20526_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6943_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_11), .I3(ootx_shift_registers_1_12), 
            .O(n11053));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6943_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_1942_24_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n22749), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6942_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_10), .I3(ootx_shift_registers_1_11), 
            .O(n11052));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6942_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7152_3_lut_4_lut (.I0(n1004), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_241), .O(n11262));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7152_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i92_2_lut (.I0(n60_adj_2038), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i92_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mod_155_add_1808_24_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n22698), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_355_21 (.CI(n22293), .I0(\counter_from_last_rise[19] ), 
            .I1(GND_net), .CO(n22294));
    SB_LUT4 i7743_3_lut_4_lut (.I0(n1002), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1193), .O(n11853));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7743_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6941_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_9), .I3(ootx_shift_registers_1_10), 
            .O(n11051));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6941_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7151_3_lut_4_lut (.I0(n1002), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_240), .O(n11261));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7151_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7563_3_lut_4_lut (.I0(n642), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1373), .O(n11673));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i359_360_adj_863 (.Q(ootx_payloads_0_27), .C(clock_c), .D(n10982));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i13_4_lut_adj_864 (.I0(n2208), .I1(n2197), .I2(n2201), .I3(n2202), 
            .O(n31_adj_2238));
    defparam i13_4_lut_adj_864.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1540_19 (.CI(n22603), .I0(n2196), .I1(n2225), 
            .CO(n22604));
    SB_LUT4 mod_155_add_2143_4_lut (.I0(n3112_c), .I1(n3112_c), .I2(n3116), 
            .I3(n22813), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7007_3_lut_4_lut (.I0(n714), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_96), .O(n11117));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7007_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7599_3_lut_4_lut (.I0(n714), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1337), .O(n11709));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6971_3_lut_4_lut (.I0(n642), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_60), .O(n11081));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6971_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_865 (.I0(n2851[10]), .I1(n2212), .I2(n2211), 
            .I3(n2210), .O(n22947));
    defparam i3_4_lut_adj_865.LUT_INIT = 16'hfffe;
    SB_DFF i389_390_adj_866 (.Q(ootx_payloads_0_37), .C(clock_c), .D(n10981));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 mod_155_add_1071_13_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n22478), .O(n1601_adj_2150)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_2143_4 (.CI(n22813), .I0(n3112_c), .I1(n3116), 
            .CO(n22814));
    SB_LUT4 i4_2_lut_adj_867 (.I0(n2192), .I1(n2200), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_2239));
    defparam i4_2_lut_adj_867.LUT_INIT = 16'heeee;
    SB_LUT4 Mux_31_i1_3_lut_adj_868 (.I0(bit_counters_0_5), .I1(bit_counters_1_5), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[5]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_31_i1_3_lut_adj_868.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_869 (.I0(n2203), .I1(n2206), .I2(n2199), .I3(n2205), 
            .O(n30_adj_2240));
    defparam i12_4_lut_adj_869.LUT_INIT = 16'hfffe;
    SB_CARRY mod_155_add_1071_13 (.CI(n22478), .I0(n1502), .I1(n1532), 
            .CO(n22479));
    SB_DFF i383_384_adj_870 (.Q(ootx_payloads_0_35), .C(clock_c), .D(n10980));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_CARRY mod_155_add_2076_2 (.CI(VCC_net), .I0(n2851[2]), .I1(n25183), 
            .CO(n22783));
    SB_LUT4 i6991_3_lut_4_lut (.I0(n682), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_80), .O(n11101));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i6991_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7583_3_lut_4_lut (.I0(n682), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1353), .O(n11693));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7583_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7014_3_lut_4_lut (.I0(n728), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_103), .O(n11124));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7014_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 Mux_30_i1_3_lut_adj_871 (.I0(bit_counters_0_6), .I1(bit_counters_1_6), 
            .I2(\lighthouse[0] ), .I3(GND_net), .O(n2849[6]));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(167[24:34])
    defparam Mux_30_i1_3_lut_adj_871.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_from_nskip_rise_640_add_4_8_lut (.I0(n6359), .I1(n2280), 
            .I2(counter_from_nskip_rise[6]), .I3(n22356), .O(n91[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_from_nskip_rise_640_add_4_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mod_155_add_1942_24 (.CI(n22749), .I0(n2791), .I1(n2819), 
            .CO(n22750));
    SB_LUT4 i16_4_lut_adj_872 (.I0(n31_adj_2238), .I1(n2195), .I2(n28_adj_2237), 
            .I3(n2193), .O(n34_adj_2241));
    defparam i16_4_lut_adj_872.LUT_INIT = 16'hfffe;
    SB_LUT4 i6940_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_8), .I3(ootx_shift_registers_1_9), 
            .O(n11050));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6940_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7606_3_lut_4_lut (.I0(n728), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1330), .O(n11716));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7606_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_3_lut_adj_873 (.I0(n2196), .I1(n22947), .I2(n2209), .I3(GND_net), 
            .O(n21_adj_2242));
    defparam i3_3_lut_adj_873.LUT_INIT = 16'heaea;
    SB_DFFESR sync__i0 (.Q(sync[0]), .C(clock_c), .E(n2282), .D(n112), 
            .R(n18844));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 i6939_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_7), .I3(ootx_shift_registers_1_8), 
            .O(n11049));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6939_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mod_155_add_1540_18_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n22602), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6938_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_6), .I3(ootx_shift_registers_1_7), 
            .O(n11048));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6938_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY mod_155_add_1808_24 (.CI(n22698), .I0(n2591), .I1(n2621), 
            .CO(n22699));
    SB_LUT4 i6937_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_5), .I3(ootx_shift_registers_1_6), 
            .O(n11047));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6937_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i17_4_lut_adj_874 (.I0(n21_adj_2242), .I1(n34_adj_2241), .I2(n30_adj_2240), 
            .I3(n22_adj_2239), .O(n2225));
    defparam i17_4_lut_adj_874.LUT_INIT = 16'hfffe;
    SB_DFFER led_i0_i8 (.Q(led_c_7), .C(clock_c), .E(n23741), .D(n4731), 
            .R(reset_c));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(82[4] 343[11])
    SB_LUT4 mod_155_add_1071_12_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n22477), .O(n1602_adj_2154)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_155_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_155_add_1540_18 (.CI(n22602), .I0(n2197), .I1(n2225), 
            .CO(n22603));
    SB_LUT4 i6936_3_lut_4_lut (.I0(ootx_shift_registers_N_1748), .I1(\lighthouse[0] ), 
            .I2(ootx_shift_registers_1_4), .I3(ootx_shift_registers_1_5), 
            .O(n11046));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(92[41:42])
    defparam i6936_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut (.I0(n40_adj_2049), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n88_adj_1877));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i88_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut (.I0(n40_adj_2049), .I1(\ootx_payloads_N_1699[4] ), 
            .I2(\ootx_payloads_N_1699[5] ), .I3(GND_net), .O(n87));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i87_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i650_651_adj_875 (.Q(ootx_payloads_0_124), .C(clock_c), .D(n11145));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(44[9:22])
    SB_LUT4 i7013_3_lut_4_lut (.I0(n726), .I1(\lighthouse[0] ), .I2(data), 
            .I3(ootx_payloads_0_102), .O(n11123));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7605_3_lut_4_lut (.I0(n726), .I1(\lighthouse[0] ), .I2(data), 
            .I3(n1331), .O(n11715));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam i7605_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i170_2_lut_3_lut (.I0(n41_adj_1946), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n170_adj_2042));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i170_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i169_2_lut_3_lut (.I0(n41_adj_1946), .I1(\ootx_payloads_N_1699[5] ), 
            .I2(\ootx_payloads_N_1699[6] ), .I3(GND_net), .O(n169));   // ../../roboy_control/src/roboy_plexus/roboy_de10_nano_soc/ip/roboy_fpga_code/lighthouse_tracking/lighthouse_ootx_decoder.vhdl(148[37:62])
    defparam EnabledDecoder_2_i169_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_CARRY counter_from_nskip_rise_640_add_4_8 (.CI(n22356), .I0(n2280), 
            .I1(counter_from_nskip_rise[6]), .CO(n22357));
    SB_CARRY add_154_21 (.CI(n22262), .I0(n2849[19]), .I1(GND_net), .CO(n22263));
    
endmodule
